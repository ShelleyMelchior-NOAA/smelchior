<!DOCTYPE html PUBLIC "-//w3c//dtd html 4.0 transitional//en">
<html>
<head>

  
  <meta http-equiv="Content-Type" content="text/html; charset=iso-8859-1">

  
  <meta name="Generator" content="WordPerfect 9">

  
  <meta name="GENERATOR" content="Mozilla/4.7 [en] (Win98; U) [Netscape]">

  
  <meta name="Author" content="Dennis Keyser">

  
  <title>CODE TABLE FOR INPUT REPORT TYPES</title>
</head>


<body alink="#ff0000" bgcolor="#ffffff" link="#0000ff" text="#000000" vlink="#551a8b">

&nbsp;
<br>

Table 6.&nbsp; Code table for input report types (last revised
2/12/2018)<span style="font-style: italic;"> (should be&nbsp;up-to-date)</span>.
<br>

&nbsp;
<table style="width: 100%;" border="1">

  <tbody>

    <tr valign="top">

      <td>Report Type</td>

      <td>Definition</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 11</td>

      <td>Fixed land RAOB and PIBAL by block and station number</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 12</td>

      <td>Fixed land RAOB and PIBAL by call letters</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 13</td>

      <td>Mobile land RAOB (including CLAS soundings)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 22</td>

      <td>Ship RAOB with name</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 23</td>

      <td>Ship RAOB without name (report id set to "SHIP")</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 31</td>

      <td>Reconnaissance aircraft or dropwinsonde</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 41&nbsp;</td>

      <td>Aircraft flight-level (all types)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 61</td>

      <td>Satellite soundings/retrievals/radiances</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 63</td>

      <td>Satellite-derived winds</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 65</td>

      <td>SSM/I total precipitable water (ocean) product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 66</td>

      <td>SSM/I rain rate product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 68</td>

      <td>SSM/I brightness temperatures</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 69</td>

      <td>SSM/I cloud water (ocean) product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 71</td>

      <td>NOAA Profiler Network (NPN) Profiler winds</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 72</td>

      <td>NEXRAD Vertical Azimuth Display (VAD) winds &nbsp;(from both Radar Coded Message and&nbsp;from Level 2 decoder)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 73</td>

      <td>Wind profiler originating in PIBAL bulletins (tropical
and European)</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp; &nbsp;74</td>

      <td>GPS-IPW (Integrated Precipitable Water)</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp; &nbsp;75</td>

      <td>Multi-Agency Profiler (MAP) Profiler and&nbsp;acoustic
sounder (SODAR) winds</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp; &nbsp;76</td>

      <td>Japanese Meteorological Agency (JMA) profiler winds</td>

    </tr>

    <tr>

      <td style="vertical-align: top;">&nbsp; &nbsp; &nbsp; &nbsp;
&nbsp;77</td>

      <td>NOAA Profiler Network (NPN) or Multi-Agency Profiler (MAP)
RASS temperatures</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 511</td>

      <td>Land surface (fixed) by block and station number (synoptic, both
unrestricted &amp; restricted WMO Res. 40)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 512</td>

      <td>Land surface (fixed) by call letters (METAR)</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp;514</td>

      <td>Mobile land surface (synoptic)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 522</td>

      <td>Ship with name</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 523</td>

      <td>Ship without name (report id set to "SHIP")</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 531</td>

      <td>C-MAN platform</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 532</td>

      <td>Tide gauge report</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp;534</td>

      <td>Coast&nbsp;Guard tide gauge report</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp;540</td>

      <td>Mesonet surface</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 551</td>

      <td>Sea-level pressure bogus</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 561</td>

      <td>Buoys arriving in TAC WMO FM13 format (fixed)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 562</td>

      <td>Buoys arriving in TAC WMO FM18 format (fixed or drifting)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 563</td>

      <td>Buoys arriving in BUFR format (fixed)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 564</td>

      <td>Buoys arriving in BUFR format (drifting)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 571</td>

      <td>SSM/I wind speed (ocean) product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 573</td>

      <td>SSM/I soil moisture product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 574</td>

      <td>SSM/I snow depth product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 575</td>

      <td>SSM/I additional products (surface tag, ice concentration,
ice age, ice edge, calculated surface type)</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 576</td>

      <td>SSM/I surface (skin) temperature product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 577</td>

      <td>SSM/I sea surface temperature product</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 581</td>

      <td>ERS scatterometer winds</td>

    </tr>

    <tr valign="top">

      <td>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;&nbsp; 582</td>

      <td>QuikSCAT scatterometer winds</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp;583</td>

      <td>WindSAT scatterometer winds (Navy- or NESDIS- produced)</td>

    </tr>

    <tr>

      <td>&nbsp; &nbsp; &nbsp; &nbsp;584</td>

      <td>ASCAT scatterometer winds</td>

    </tr>

  
  </tbody>
</table>

<br clear="all">

<br>

<br>

</body>
</html>

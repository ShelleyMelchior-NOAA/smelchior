<?xml version='1.0' encoding='UTF-8'?>
<kml xmlns="http://www.opengis.net/kml/2.2">
<Document>
<name>rtmamoist_aws_plot.kml</name>
<open>1</open>
<Style id='zero'>
<IconStyle>
<color>FFFFFFFF</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='ten'>
<IconStyle>
<color>FFFFFF00</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle2.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='twenty'>
<IconStyle>
<color>FFFF0000</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle3.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='thirty'>
<IconStyle>
<color>FF00FF00</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle4.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='fourty'>
<IconStyle>
<color>FF008000</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle5.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='fifty'>
<IconStyle>
<color>FF00FFFF</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle6.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='sixty'>
<IconStyle>
<color>FF008080</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle7.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='seventy'>
<IconStyle>
<color>FF0000FF</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle8.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='eighty'>
<IconStyle>
<color>FF000080</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle9.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='ninety'>
<IconStyle>
<color>FF800080</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle10.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Style id='hundred'>
<IconStyle>
<color>FFFF00FF</color>
<scale>1.5</scale>
<Icon>
<href>http://www.emc.ncep.noaa.gov/mmb/obsdumpmonitor/icon/placemark_circle11.png</href>
</Icon>
</IconStyle>
<LabelStyle>
<scale>1.5</scale>
</LabelStyle>
</Style>
<Folder name='0 AWS'>
<Placemark>
<name>23.5 N, -70.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-70.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -75.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-75.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 29 non-AWS obs</description>
<Point>
<coordinates>-81.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1 non-AWS obs</description>
<Point>
<coordinates>-82.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 9 non-AWS obs</description>
<Point>
<coordinates>-98.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 6 non-AWS obs</description>
<Point>
<coordinates>-99.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-103.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 26 non-AWS obs</description>
<Point>
<coordinates>-106.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>23.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 80 non-AWS obs</description>
<Point>
<coordinates>-109.5,23.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>24.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-80.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>24.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 263 non-AWS obs</description>
<Point>
<coordinates>-81.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>24.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 9 non-AWS obs</description>
<Point>
<coordinates>-104.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>24.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 2 non-AWS obs</description>
<Point>
<coordinates>-107.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>24.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 16 non-AWS obs</description>
<Point>
<coordinates>-110.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>25.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1 non-AWS obs</description>
<Point>
<coordinates>-103.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>25.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 2 non-AWS obs</description>
<Point>
<coordinates>-105.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>25.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1 non-AWS obs</description>
<Point>
<coordinates>-109.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>25.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-111.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 20 non-AWS obs</description>
<Point>
<coordinates>-78.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -85.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-85.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -96.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-96.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 29 non-AWS obs</description>
<Point>
<coordinates>-99.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-101.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-108.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 13 non-AWS obs</description>
<Point>
<coordinates>-111.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-71.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 80 non-AWS obs</description>
<Point>
<coordinates>-90.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-95.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 106 non-AWS obs</description>
<Point>
<coordinates>-98.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1 non-AWS obs</description>
<Point>
<coordinates>-109.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-110.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-112.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-78.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-84.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 73 non-AWS obs</description>
<Point>
<coordinates>-88.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -89.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 171 non-AWS obs</description>
<Point>
<coordinates>-89.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 16 non-AWS obs</description>
<Point>
<coordinates>-90.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-98.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 30 non-AWS obs</description>
<Point>
<coordinates>-99.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-100.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1 non-AWS obs</description>
<Point>
<coordinates>-106.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 7 non-AWS obs</description>
<Point>
<coordinates>-117.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 169 non-AWS obs</description>
<Point>
<coordinates>-83.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-84.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -85.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-85.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-88.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-92.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-103.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 7 non-AWS obs</description>
<Point>
<coordinates>-104.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-110.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 231 non-AWS obs</description>
<Point>
<coordinates>-83.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -85.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 233 non-AWS obs</description>
<Point>
<coordinates>-85.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 44 non-AWS obs</description>
<Point>
<coordinates>-101.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-102.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-103.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-107.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-69.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-80.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 264 non-AWS obs</description>
<Point>
<coordinates>-81.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 140 non-AWS obs</description>
<Point>
<coordinates>-82.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 61 non-AWS obs</description>
<Point>
<coordinates>-83.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 43 non-AWS obs</description>
<Point>
<coordinates>-84.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -87.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-87.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 102 non-AWS obs</description>
<Point>
<coordinates>-90.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 139 non-AWS obs</description>
<Point>
<coordinates>-93.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 438 non-AWS obs</description>
<Point>
<coordinates>-98.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 219 non-AWS obs</description>
<Point>
<coordinates>-99.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-101.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-103.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-105.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-81.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-82.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 200 non-AWS obs</description>
<Point>
<coordinates>-83.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 161 non-AWS obs</description>
<Point>
<coordinates>-84.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-91.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 972 non-AWS obs</description>
<Point>
<coordinates>-100.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-101.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 167 non-AWS obs</description>
<Point>
<coordinates>-102.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 212 non-AWS obs</description>
<Point>
<coordinates>-105.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 167 non-AWS obs</description>
<Point>
<coordinates>-109.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-112.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 949 non-AWS obs</description>
<Point>
<coordinates>-114.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-115.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -77.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-77.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 241 non-AWS obs</description>
<Point>
<coordinates>-78.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 274 non-AWS obs</description>
<Point>
<coordinates>-80.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 143 non-AWS obs</description>
<Point>
<coordinates>-82.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 154 non-AWS obs</description>
<Point>
<coordinates>-88.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -89.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 30 non-AWS obs</description>
<Point>
<coordinates>-89.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 76 non-AWS obs</description>
<Point>
<coordinates>-90.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 117 non-AWS obs</description>
<Point>
<coordinates>-99.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-100.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 175 non-AWS obs</description>
<Point>
<coordinates>-102.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-103.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-108.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-109.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-110.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-113.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 56 non-AWS obs</description>
<Point>
<coordinates>-114.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-115.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 273 non-AWS obs</description>
<Point>
<coordinates>-118.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 41 non-AWS obs</description>
<Point>
<coordinates>-119.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-120.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-72.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -79.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 302 non-AWS obs</description>
<Point>
<coordinates>-79.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 198 non-AWS obs</description>
<Point>
<coordinates>-95.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 369 non-AWS obs</description>
<Point>
<coordinates>-97.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 188 non-AWS obs</description>
<Point>
<coordinates>-99.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-100.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 120 non-AWS obs</description>
<Point>
<coordinates>-103.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 20 non-AWS obs</description>
<Point>
<coordinates>-104.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-108.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 719 non-AWS obs</description>
<Point>
<coordinates>-109.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 148 non-AWS obs</description>
<Point>
<coordinates>-110.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 336 non-AWS obs</description>
<Point>
<coordinates>-111.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 59 non-AWS obs</description>
<Point>
<coordinates>-113.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 181 non-AWS obs</description>
<Point>
<coordinates>-120.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -75.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 62 non-AWS obs</description>
<Point>
<coordinates>-75.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -76.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-76.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 289 non-AWS obs</description>
<Point>
<coordinates>-98.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 146 non-AWS obs</description>
<Point>
<coordinates>-99.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 132 non-AWS obs</description>
<Point>
<coordinates>-100.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-101.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-102.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 58 non-AWS obs</description>
<Point>
<coordinates>-110.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 201 non-AWS obs</description>
<Point>
<coordinates>-111.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-112.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 155 non-AWS obs</description>
<Point>
<coordinates>-113.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-115.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-116.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 168 non-AWS obs</description>
<Point>
<coordinates>-117.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 448 non-AWS obs</description>
<Point>
<coordinates>-118.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 256 non-AWS obs</description>
<Point>
<coordinates>-120.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-121.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-74.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 30 non-AWS obs</description>
<Point>
<coordinates>-91.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 109 non-AWS obs</description>
<Point>
<coordinates>-92.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 172 non-AWS obs</description>
<Point>
<coordinates>-93.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 435 non-AWS obs</description>
<Point>
<coordinates>-97.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 296 non-AWS obs</description>
<Point>
<coordinates>-99.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 564 non-AWS obs</description>
<Point>
<coordinates>-101.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-102.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-103.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-106.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 19 non-AWS obs</description>
<Point>
<coordinates>-109.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 191 non-AWS obs</description>
<Point>
<coordinates>-111.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 67 non-AWS obs</description>
<Point>
<coordinates>-112.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-113.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 92 non-AWS obs</description>
<Point>
<coordinates>-120.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 149 non-AWS obs</description>
<Point>
<coordinates>-92.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-106.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-108.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 504 non-AWS obs</description>
<Point>
<coordinates>-116.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 2 non-AWS obs</description>
<Point>
<coordinates>-117.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 499 non-AWS obs</description>
<Point>
<coordinates>-119.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-80.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 113 non-AWS obs</description>
<Point>
<coordinates>-81.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 117 non-AWS obs</description>
<Point>
<coordinates>-102.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 201 non-AWS obs</description>
<Point>
<coordinates>-107.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 167 non-AWS obs</description>
<Point>
<coordinates>-108.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-109.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 67 non-AWS obs</description>
<Point>
<coordinates>-110.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 14 non-AWS obs</description>
<Point>
<coordinates>-116.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 92 non-AWS obs</description>
<Point>
<coordinates>-123.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 82 non-AWS obs</description>
<Point>
<coordinates>-72.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 74 non-AWS obs</description>
<Point>
<coordinates>-91.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-92.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 226 non-AWS obs</description>
<Point>
<coordinates>-107.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-109.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 727 non-AWS obs</description>
<Point>
<coordinates>-112.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-113.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 97 non-AWS obs</description>
<Point>
<coordinates>-116.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 190 non-AWS obs</description>
<Point>
<coordinates>-117.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 49 non-AWS obs</description>
<Point>
<coordinates>-118.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 166 non-AWS obs</description>
<Point>
<coordinates>-120.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 303 non-AWS obs</description>
<Point>
<coordinates>-121.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 311 non-AWS obs</description>
<Point>
<coordinates>-122.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 223 non-AWS obs</description>
<Point>
<coordinates>-123.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 134 non-AWS obs</description>
<Point>
<coordinates>-90.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 150 non-AWS obs</description>
<Point>
<coordinates>-92.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -94.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 136 non-AWS obs</description>
<Point>
<coordinates>-94.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 143 non-AWS obs</description>
<Point>
<coordinates>-98.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-103.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 139 non-AWS obs</description>
<Point>
<coordinates>-107.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 52 non-AWS obs</description>
<Point>
<coordinates>-108.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 444 non-AWS obs</description>
<Point>
<coordinates>-113.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-118.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-119.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 223 non-AWS obs</description>
<Point>
<coordinates>-120.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 195 non-AWS obs</description>
<Point>
<coordinates>-121.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 666 non-AWS obs</description>
<Point>
<coordinates>-122.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 157 non-AWS obs</description>
<Point>
<coordinates>-123.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -124.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-124.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 76 non-AWS obs</description>
<Point>
<coordinates>-69.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 186 non-AWS obs</description>
<Point>
<coordinates>-90.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 457 non-AWS obs</description>
<Point>
<coordinates>-95.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-98.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-99.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-105.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 136 non-AWS obs</description>
<Point>
<coordinates>-106.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-107.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-113.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-115.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-116.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-118.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-119.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 214 non-AWS obs</description>
<Point>
<coordinates>-120.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 164 non-AWS obs</description>
<Point>
<coordinates>-121.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 260 non-AWS obs</description>
<Point>
<coordinates>-123.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 113 non-AWS obs</description>
<Point>
<coordinates>-74.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 51 non-AWS obs</description>
<Point>
<coordinates>-80.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-81.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -96.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 268 non-AWS obs</description>
<Point>
<coordinates>-96.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 14 non-AWS obs</description>
<Point>
<coordinates>-99.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 77 non-AWS obs</description>
<Point>
<coordinates>-100.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 65 non-AWS obs</description>
<Point>
<coordinates>-101.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-103.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-104.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-105.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-106.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 55 non-AWS obs</description>
<Point>
<coordinates>-107.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-108.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 73 non-AWS obs</description>
<Point>
<coordinates>-110.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-111.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 296 non-AWS obs</description>
<Point>
<coordinates>-112.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 355 non-AWS obs</description>
<Point>
<coordinates>-113.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 93 non-AWS obs</description>
<Point>
<coordinates>-115.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-116.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 9 non-AWS obs</description>
<Point>
<coordinates>-117.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-119.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 87 non-AWS obs</description>
<Point>
<coordinates>-120.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 190 non-AWS obs</description>
<Point>
<coordinates>-121.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 249 non-AWS obs</description>
<Point>
<coordinates>-122.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 266 non-AWS obs</description>
<Point>
<coordinates>-123.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -124.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 11 non-AWS obs</description>
<Point>
<coordinates>-124.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-66.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-68.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 146 non-AWS obs</description>
<Point>
<coordinates>-80.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-81.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 217 non-AWS obs</description>
<Point>
<coordinates>-82.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -94.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 171 non-AWS obs</description>
<Point>
<coordinates>-94.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -96.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 418 non-AWS obs</description>
<Point>
<coordinates>-96.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 92 non-AWS obs</description>
<Point>
<coordinates>-98.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-99.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-100.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-101.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-102.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-105.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-106.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-107.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-108.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-109.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 307 non-AWS obs</description>
<Point>
<coordinates>-110.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 202 non-AWS obs</description>
<Point>
<coordinates>-111.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 2910 non-AWS obs</description>
<Point>
<coordinates>-112.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 138 non-AWS obs</description>
<Point>
<coordinates>-115.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-118.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 26 non-AWS obs</description>
<Point>
<coordinates>-119.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 133 non-AWS obs</description>
<Point>
<coordinates>-121.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 101 non-AWS obs</description>
<Point>
<coordinates>-122.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 168 non-AWS obs</description>
<Point>
<coordinates>-123.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -124.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-124.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-66.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -67.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-67.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 475 non-AWS obs</description>
<Point>
<coordinates>-68.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 290 non-AWS obs</description>
<Point>
<coordinates>-69.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -70.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 186 non-AWS obs</description>
<Point>
<coordinates>-70.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -73.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 377 non-AWS obs</description>
<Point>
<coordinates>-73.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 184 non-AWS obs</description>
<Point>
<coordinates>-74.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -76.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 140 non-AWS obs</description>
<Point>
<coordinates>-76.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -77.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-77.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-78.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -79.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1087 non-AWS obs</description>
<Point>
<coordinates>-79.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-81.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-82.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-83.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 213 non-AWS obs</description>
<Point>
<coordinates>-84.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -86.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 82 non-AWS obs</description>
<Point>
<coordinates>-86.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -96.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 350 non-AWS obs</description>
<Point>
<coordinates>-96.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 191 non-AWS obs</description>
<Point>
<coordinates>-97.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 114 non-AWS obs</description>
<Point>
<coordinates>-98.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-99.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 144 non-AWS obs</description>
<Point>
<coordinates>-100.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-101.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-105.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 135 non-AWS obs</description>
<Point>
<coordinates>-108.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-109.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-110.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 92 non-AWS obs</description>
<Point>
<coordinates>-111.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 475 non-AWS obs</description>
<Point>
<coordinates>-112.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 107 non-AWS obs</description>
<Point>
<coordinates>-113.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 137 non-AWS obs</description>
<Point>
<coordinates>-114.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-115.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 153 non-AWS obs</description>
<Point>
<coordinates>-117.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 55 non-AWS obs</description>
<Point>
<coordinates>-118.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-120.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 155 non-AWS obs</description>
<Point>
<coordinates>-66.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -67.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-67.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-68.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-69.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-71.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 54 non-AWS obs</description>
<Point>
<coordinates>-72.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -73.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 305 non-AWS obs</description>
<Point>
<coordinates>-73.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 51 non-AWS obs</description>
<Point>
<coordinates>-74.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -75.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-75.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -76.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-76.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -77.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 65 non-AWS obs</description>
<Point>
<coordinates>-77.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-78.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -79.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-79.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-80.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 25 non-AWS obs</description>
<Point>
<coordinates>-81.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-82.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-83.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -85.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 126 non-AWS obs</description>
<Point>
<coordinates>-85.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -86.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 65 non-AWS obs</description>
<Point>
<coordinates>-86.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 120 non-AWS obs</description>
<Point>
<coordinates>-90.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-97.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-98.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-99.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-101.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-102.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-103.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 25 non-AWS obs</description>
<Point>
<coordinates>-104.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-107.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-108.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-109.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 152 non-AWS obs</description>
<Point>
<coordinates>-111.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 78 non-AWS obs</description>
<Point>
<coordinates>-112.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 182 non-AWS obs</description>
<Point>
<coordinates>-113.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-114.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 51 non-AWS obs</description>
<Point>
<coordinates>-115.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 128 non-AWS obs</description>
<Point>
<coordinates>-116.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 203 non-AWS obs</description>
<Point>
<coordinates>-117.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 225 non-AWS obs</description>
<Point>
<coordinates>-119.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -124.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-124.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -67.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 108 non-AWS obs</description>
<Point>
<coordinates>-67.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 135 non-AWS obs</description>
<Point>
<coordinates>-68.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-69.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -70.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-70.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 133 non-AWS obs</description>
<Point>
<coordinates>-71.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-72.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-74.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -75.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 3 non-AWS obs</description>
<Point>
<coordinates>-75.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-80.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 20 non-AWS obs</description>
<Point>
<coordinates>-81.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-83.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 158 non-AWS obs</description>
<Point>
<coordinates>-84.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -85.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-85.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -86.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 107 non-AWS obs</description>
<Point>
<coordinates>-86.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -87.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 131 non-AWS obs</description>
<Point>
<coordinates>-87.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 68 non-AWS obs</description>
<Point>
<coordinates>-88.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -89.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-89.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 187 non-AWS obs</description>
<Point>
<coordinates>-90.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-97.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-99.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-100.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-101.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-102.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-103.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-104.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 76 non-AWS obs</description>
<Point>
<coordinates>-105.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 6 non-AWS obs</description>
<Point>
<coordinates>-106.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 132 non-AWS obs</description>
<Point>
<coordinates>-108.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-109.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-110.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 115 non-AWS obs</description>
<Point>
<coordinates>-111.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 133 non-AWS obs</description>
<Point>
<coordinates>-112.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 139 non-AWS obs</description>
<Point>
<coordinates>-113.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 133 non-AWS obs</description>
<Point>
<coordinates>-114.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 44 non-AWS obs</description>
<Point>
<coordinates>-115.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 195 non-AWS obs</description>
<Point>
<coordinates>-116.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 191 non-AWS obs</description>
<Point>
<coordinates>-118.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 101 non-AWS obs</description>
<Point>
<coordinates>-120.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 19 non-AWS obs</description>
<Point>
<coordinates>-66.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -67.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-67.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-69.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -70.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 59 non-AWS obs</description>
<Point>
<coordinates>-70.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 44 non-AWS obs</description>
<Point>
<coordinates>-71.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-72.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-74.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -79.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 73 non-AWS obs</description>
<Point>
<coordinates>-79.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -83.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 19 non-AWS obs</description>
<Point>
<coordinates>-83.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-84.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -87.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-87.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-88.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -89.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-89.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-90.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 164 non-AWS obs</description>
<Point>
<coordinates>-91.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 228 non-AWS obs</description>
<Point>
<coordinates>-92.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-93.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-95.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 136 non-AWS obs</description>
<Point>
<coordinates>-97.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-98.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -99.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-99.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -100.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-100.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 41 non-AWS obs</description>
<Point>
<coordinates>-102.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-103.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 97 non-AWS obs</description>
<Point>
<coordinates>-104.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-105.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 53 non-AWS obs</description>
<Point>
<coordinates>-106.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-107.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 87 non-AWS obs</description>
<Point>
<coordinates>-108.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-109.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 67 non-AWS obs</description>
<Point>
<coordinates>-110.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-111.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-113.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 219 non-AWS obs</description>
<Point>
<coordinates>-114.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 193 non-AWS obs</description>
<Point>
<coordinates>-115.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -67.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 16 non-AWS obs</description>
<Point>
<coordinates>-67.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 30 non-AWS obs</description>
<Point>
<coordinates>-68.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -69.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-69.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -70.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 44 non-AWS obs</description>
<Point>
<coordinates>-70.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-71.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -72.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 54 non-AWS obs</description>
<Point>
<coordinates>-72.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -77.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 56 non-AWS obs</description>
<Point>
<coordinates>-77.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-78.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -79.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 37 non-AWS obs</description>
<Point>
<coordinates>-79.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -81.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 146 non-AWS obs</description>
<Point>
<coordinates>-81.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -86.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-86.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -87.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-87.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-90.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 3 non-AWS obs</description>
<Point>
<coordinates>-91.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 115 non-AWS obs</description>
<Point>
<coordinates>-92.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 157 non-AWS obs</description>
<Point>
<coordinates>-93.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -94.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 117 non-AWS obs</description>
<Point>
<coordinates>-94.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 141 non-AWS obs</description>
<Point>
<coordinates>-95.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -96.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-96.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-97.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -98.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-98.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -101.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-101.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 51 non-AWS obs</description>
<Point>
<coordinates>-102.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 60 non-AWS obs</description>
<Point>
<coordinates>-104.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 77 non-AWS obs</description>
<Point>
<coordinates>-105.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 142 non-AWS obs</description>
<Point>
<coordinates>-106.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 77 non-AWS obs</description>
<Point>
<coordinates>-107.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-108.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-109.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 29 non-AWS obs</description>
<Point>
<coordinates>-110.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-111.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-112.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -113.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-113.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-115.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 61 non-AWS obs</description>
<Point>
<coordinates>-120.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-66.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -68.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 44 non-AWS obs</description>
<Point>
<coordinates>-68.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -71.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-71.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -74.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-74.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -77.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-77.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -82.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 55 non-AWS obs</description>
<Point>
<coordinates>-82.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-84.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -86.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-86.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -88.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-88.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 17 non-AWS obs</description>
<Point>
<coordinates>-90.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -92.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-92.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-93.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -94.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 87 non-AWS obs</description>
<Point>
<coordinates>-94.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-102.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-103.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 35 non-AWS obs</description>
<Point>
<coordinates>-105.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-107.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -108.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-108.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-109.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 35 non-AWS obs</description>
<Point>
<coordinates>-114.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-115.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 55 non-AWS obs</description>
<Point>
<coordinates>-117.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 175 non-AWS obs</description>
<Point>
<coordinates>-119.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 43 non-AWS obs</description>
<Point>
<coordinates>-120.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 60 non-AWS obs</description>
<Point>
<coordinates>-121.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 274 non-AWS obs</description>
<Point>
<coordinates>-122.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -124.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 312 non-AWS obs</description>
<Point>
<coordinates>-124.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -125.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-125.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -126.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 36 non-AWS obs</description>
<Point>
<coordinates>-126.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -66.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-66.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -91.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-91.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 11 non-AWS obs</description>
<Point>
<coordinates>-93.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 15 non-AWS obs</description>
<Point>
<coordinates>-95.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-102.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -103.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-103.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 86 non-AWS obs</description>
<Point>
<coordinates>-104.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 42 non-AWS obs</description>
<Point>
<coordinates>-105.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 213 non-AWS obs</description>
<Point>
<coordinates>-107.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-109.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -114.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-114.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -117.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 26 non-AWS obs</description>
<Point>
<coordinates>-117.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -118.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 14 non-AWS obs</description>
<Point>
<coordinates>-118.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -119.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-119.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -120.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 75 non-AWS obs</description>
<Point>
<coordinates>-120.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 176 non-AWS obs</description>
<Point>
<coordinates>-121.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -122.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 1499 non-AWS obs</description>
<Point>
<coordinates>-122.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -123.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 54 non-AWS obs</description>
<Point>
<coordinates>-123.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -127.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-127.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -76.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-76.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -78.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 9 non-AWS obs</description>
<Point>
<coordinates>-78.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -80.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 60 non-AWS obs</description>
<Point>
<coordinates>-80.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -90.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 83 non-AWS obs</description>
<Point>
<coordinates>-90.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -93.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-93.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -95.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 14 non-AWS obs</description>
<Point>
<coordinates>-95.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -102.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-102.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -104.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-104.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -105.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 56 non-AWS obs</description>
<Point>
<coordinates>-105.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-106.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -107.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-107.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-109.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -115.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 56 non-AWS obs</description>
<Point>
<coordinates>-115.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-116.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-121.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -127.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 33 non-AWS obs</description>
<Point>
<coordinates>-127.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -87.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-87.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -97.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-97.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -106.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-106.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 68 non-AWS obs</description>
<Point>
<coordinates>-110.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 131 non-AWS obs</description>
<Point>
<coordinates>-111.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -112.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 189 non-AWS obs</description>
<Point>
<coordinates>-112.5,52.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -84.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-84.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -94.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 15 non-AWS obs</description>
<Point>
<coordinates>-94.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -109.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 15 non-AWS obs</description>
<Point>
<coordinates>-109.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -110.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 18 non-AWS obs</description>
<Point>
<coordinates>-110.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -111.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 52 non-AWS obs</description>
<Point>
<coordinates>-111.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -116.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 14 non-AWS obs</description>
<Point>
<coordinates>-116.5,53.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>53.5 N, -121.5 W</name>
<styleUrl>#zero</styleUrl>
<description>0 AWS obs, 13 non-AWS obs</description>
<Point>
<coordinates>-121.5,53.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='1-10% AWS'>
<Placemark>
<name>25.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>43 AWS obs, 427 non-AWS obs</description>
<Point>
<coordinates>-81.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>53 AWS obs, 1025 non-AWS obs</description>
<Point>
<coordinates>-81.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -97.5 W</name>
<styleUrl>#ten</styleUrl>
<description>14 AWS obs, 326 non-AWS obs</description>
<Point>
<coordinates>-97.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -80.5 W</name>
<styleUrl>#ten</styleUrl>
<description>54 AWS obs, 599 non-AWS obs</description>
<Point>
<coordinates>-80.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 485 non-AWS obs</description>
<Point>
<coordinates>-96.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>36 AWS obs, 521 non-AWS obs</description>
<Point>
<coordinates>-81.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -98.5 W</name>
<styleUrl>#ten</styleUrl>
<description>30 AWS obs, 2316 non-AWS obs</description>
<Point>
<coordinates>-98.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -99.5 W</name>
<styleUrl>#ten</styleUrl>
<description>32 AWS obs, 776 non-AWS obs</description>
<Point>
<coordinates>-99.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -92.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 300 non-AWS obs</description>
<Point>
<coordinates>-92.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -100.5 W</name>
<styleUrl>#ten</styleUrl>
<description>14 AWS obs, 184 non-AWS obs</description>
<Point>
<coordinates>-100.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -110.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 326 non-AWS obs</description>
<Point>
<coordinates>-110.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -80.5 W</name>
<styleUrl>#ten</styleUrl>
<description>26 AWS obs, 268 non-AWS obs</description>
<Point>
<coordinates>-80.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -86.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 165 non-AWS obs</description>
<Point>
<coordinates>-86.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -93.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 281 non-AWS obs</description>
<Point>
<coordinates>-93.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -110.5 W</name>
<styleUrl>#ten</styleUrl>
<description>32 AWS obs, 299 non-AWS obs</description>
<Point>
<coordinates>-110.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -116.5 W</name>
<styleUrl>#ten</styleUrl>
<description>40 AWS obs, 1063 non-AWS obs</description>
<Point>
<coordinates>-116.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -117.5 W</name>
<styleUrl>#ten</styleUrl>
<description>28 AWS obs, 317 non-AWS obs</description>
<Point>
<coordinates>-117.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -83.5 W</name>
<styleUrl>#ten</styleUrl>
<description>32 AWS obs, 380 non-AWS obs</description>
<Point>
<coordinates>-83.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -87.5 W</name>
<styleUrl>#ten</styleUrl>
<description>19 AWS obs, 215 non-AWS obs</description>
<Point>
<coordinates>-87.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -101.5 W</name>
<styleUrl>#ten</styleUrl>
<description>24 AWS obs, 240 non-AWS obs</description>
<Point>
<coordinates>-101.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -104.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 1086 non-AWS obs</description>
<Point>
<coordinates>-104.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -106.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 123 non-AWS obs</description>
<Point>
<coordinates>-106.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -116.5 W</name>
<styleUrl>#ten</styleUrl>
<description>54 AWS obs, 868 non-AWS obs</description>
<Point>
<coordinates>-116.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -117.5 W</name>
<styleUrl>#ten</styleUrl>
<description>120 AWS obs, 1249 non-AWS obs</description>
<Point>
<coordinates>-117.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -76.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 248 non-AWS obs</description>
<Point>
<coordinates>-76.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -77.5 W</name>
<styleUrl>#ten</styleUrl>
<description>12 AWS obs, 253 non-AWS obs</description>
<Point>
<coordinates>-77.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>6 AWS obs, 250 non-AWS obs</description>
<Point>
<coordinates>-81.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -82.5 W</name>
<styleUrl>#ten</styleUrl>
<description>7 AWS obs, 363 non-AWS obs</description>
<Point>
<coordinates>-82.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -83.5 W</name>
<styleUrl>#ten</styleUrl>
<description>26 AWS obs, 288 non-AWS obs</description>
<Point>
<coordinates>-83.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -85.5 W</name>
<styleUrl>#ten</styleUrl>
<description>19 AWS obs, 694 non-AWS obs</description>
<Point>
<coordinates>-85.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -94.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 156 non-AWS obs</description>
<Point>
<coordinates>-94.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 241 non-AWS obs</description>
<Point>
<coordinates>-96.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -98.5 W</name>
<styleUrl>#ten</styleUrl>
<description>32 AWS obs, 301 non-AWS obs</description>
<Point>
<coordinates>-98.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -102.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 232 non-AWS obs</description>
<Point>
<coordinates>-102.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -106.5 W</name>
<styleUrl>#ten</styleUrl>
<description>12 AWS obs, 111 non-AWS obs</description>
<Point>
<coordinates>-106.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -112.5 W</name>
<styleUrl>#ten</styleUrl>
<description>29 AWS obs, 264 non-AWS obs</description>
<Point>
<coordinates>-112.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 514 non-AWS obs</description>
<Point>
<coordinates>-119.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -77.5 W</name>
<styleUrl>#ten</styleUrl>
<description>16 AWS obs, 388 non-AWS obs</description>
<Point>
<coordinates>-77.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -83.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 394 non-AWS obs</description>
<Point>
<coordinates>-83.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -86.5 W</name>
<styleUrl>#ten</styleUrl>
<description>2 AWS obs, 199 non-AWS obs</description>
<Point>
<coordinates>-86.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -91.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 176 non-AWS obs</description>
<Point>
<coordinates>-91.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -95.5 W</name>
<styleUrl>#ten</styleUrl>
<description>26 AWS obs, 316 non-AWS obs</description>
<Point>
<coordinates>-95.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>21 AWS obs, 233 non-AWS obs</description>
<Point>
<coordinates>-96.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -97.5 W</name>
<styleUrl>#ten</styleUrl>
<description>7 AWS obs, 434 non-AWS obs</description>
<Point>
<coordinates>-97.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -107.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 104 non-AWS obs</description>
<Point>
<coordinates>-107.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>12 AWS obs, 204 non-AWS obs</description>
<Point>
<coordinates>-119.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -78.5 W</name>
<styleUrl>#ten</styleUrl>
<description>26 AWS obs, 277 non-AWS obs</description>
<Point>
<coordinates>-78.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -85.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 92 non-AWS obs</description>
<Point>
<coordinates>-85.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -87.5 W</name>
<styleUrl>#ten</styleUrl>
<description>14 AWS obs, 304 non-AWS obs</description>
<Point>
<coordinates>-87.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -89.5 W</name>
<styleUrl>#ten</styleUrl>
<description>29 AWS obs, 301 non-AWS obs</description>
<Point>
<coordinates>-89.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -98.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 186 non-AWS obs</description>
<Point>
<coordinates>-98.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -117.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 82 non-AWS obs</description>
<Point>
<coordinates>-117.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -118.5 W</name>
<styleUrl>#ten</styleUrl>
<description>7 AWS obs, 183 non-AWS obs</description>
<Point>
<coordinates>-118.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 326 non-AWS obs</description>
<Point>
<coordinates>-119.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 156 non-AWS obs</description>
<Point>
<coordinates>-81.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -105.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 116 non-AWS obs</description>
<Point>
<coordinates>-105.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -107.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 342 non-AWS obs</description>
<Point>
<coordinates>-107.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -115.5 W</name>
<styleUrl>#ten</styleUrl>
<description>7 AWS obs, 133 non-AWS obs</description>
<Point>
<coordinates>-115.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -118.5 W</name>
<styleUrl>#ten</styleUrl>
<description>13 AWS obs, 127 non-AWS obs</description>
<Point>
<coordinates>-118.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -121.5 W</name>
<styleUrl>#ten</styleUrl>
<description>67 AWS obs, 716 non-AWS obs</description>
<Point>
<coordinates>-121.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -122.5 W</name>
<styleUrl>#ten</styleUrl>
<description>77 AWS obs, 1104 non-AWS obs</description>
<Point>
<coordinates>-122.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -75.5 W</name>
<styleUrl>#ten</styleUrl>
<description>67 AWS obs, 632 non-AWS obs</description>
<Point>
<coordinates>-75.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -88.5 W</name>
<styleUrl>#ten</styleUrl>
<description>34 AWS obs, 467 non-AWS obs</description>
<Point>
<coordinates>-88.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -92.5 W</name>
<styleUrl>#ten</styleUrl>
<description>4 AWS obs, 301 non-AWS obs</description>
<Point>
<coordinates>-92.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -93.5 W</name>
<styleUrl>#ten</styleUrl>
<description>16 AWS obs, 200 non-AWS obs</description>
<Point>
<coordinates>-93.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -101.5 W</name>
<styleUrl>#ten</styleUrl>
<description>5 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-101.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -103.5 W</name>
<styleUrl>#ten</styleUrl>
<description>6 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-103.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 213 non-AWS obs</description>
<Point>
<coordinates>-119.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -120.5 W</name>
<styleUrl>#ten</styleUrl>
<description>8 AWS obs, 343 non-AWS obs</description>
<Point>
<coordinates>-120.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -122.5 W</name>
<styleUrl>#ten</styleUrl>
<description>35 AWS obs, 492 non-AWS obs</description>
<Point>
<coordinates>-122.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -81.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 247 non-AWS obs</description>
<Point>
<coordinates>-81.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -104.5 W</name>
<styleUrl>#ten</styleUrl>
<description>99 AWS obs, 1306 non-AWS obs</description>
<Point>
<coordinates>-104.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -105.5 W</name>
<styleUrl>#ten</styleUrl>
<description>47 AWS obs, 1261 non-AWS obs</description>
<Point>
<coordinates>-105.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -106.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 399 non-AWS obs</description>
<Point>
<coordinates>-106.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -88.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 392 non-AWS obs</description>
<Point>
<coordinates>-88.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -89.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 270 non-AWS obs</description>
<Point>
<coordinates>-89.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -91.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 176 non-AWS obs</description>
<Point>
<coordinates>-91.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -93.5 W</name>
<styleUrl>#ten</styleUrl>
<description>14 AWS obs, 176 non-AWS obs</description>
<Point>
<coordinates>-93.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -95.5 W</name>
<styleUrl>#ten</styleUrl>
<description>26 AWS obs, 235 non-AWS obs</description>
<Point>
<coordinates>-95.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -97.5 W</name>
<styleUrl>#ten</styleUrl>
<description>8 AWS obs, 165 non-AWS obs</description>
<Point>
<coordinates>-97.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -104.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 357 non-AWS obs</description>
<Point>
<coordinates>-104.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -105.5 W</name>
<styleUrl>#ten</styleUrl>
<description>68 AWS obs, 10954 non-AWS obs</description>
<Point>
<coordinates>-105.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -106.5 W</name>
<styleUrl>#ten</styleUrl>
<description>31 AWS obs, 375 non-AWS obs</description>
<Point>
<coordinates>-106.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -111.5 W</name>
<styleUrl>#ten</styleUrl>
<description>389 AWS obs, 4388 non-AWS obs</description>
<Point>
<coordinates>-111.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -112.5 W</name>
<styleUrl>#ten</styleUrl>
<description>31 AWS obs, 2413 non-AWS obs</description>
<Point>
<coordinates>-112.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -89.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 187 non-AWS obs</description>
<Point>
<coordinates>-89.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -91.5 W</name>
<styleUrl>#ten</styleUrl>
<description>23 AWS obs, 280 non-AWS obs</description>
<Point>
<coordinates>-91.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -92.5 W</name>
<styleUrl>#ten</styleUrl>
<description>20 AWS obs, 434 non-AWS obs</description>
<Point>
<coordinates>-92.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -93.5 W</name>
<styleUrl>#ten</styleUrl>
<description>19 AWS obs, 821 non-AWS obs</description>
<Point>
<coordinates>-93.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -94.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 319 non-AWS obs</description>
<Point>
<coordinates>-94.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>42 AWS obs, 427 non-AWS obs</description>
<Point>
<coordinates>-96.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -103.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 145 non-AWS obs</description>
<Point>
<coordinates>-103.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -111.5 W</name>
<styleUrl>#ten</styleUrl>
<description>124 AWS obs, 1445 non-AWS obs</description>
<Point>
<coordinates>-111.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -112.5 W</name>
<styleUrl>#ten</styleUrl>
<description>56 AWS obs, 593 non-AWS obs</description>
<Point>
<coordinates>-112.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -122.5 W</name>
<styleUrl>#ten</styleUrl>
<description>8 AWS obs, 454 non-AWS obs</description>
<Point>
<coordinates>-122.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -73.5 W</name>
<styleUrl>#ten</styleUrl>
<description>44 AWS obs, 442 non-AWS obs</description>
<Point>
<coordinates>-73.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -75.5 W</name>
<styleUrl>#ten</styleUrl>
<description>36 AWS obs, 376 non-AWS obs</description>
<Point>
<coordinates>-75.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -89.5 W</name>
<styleUrl>#ten</styleUrl>
<description>19 AWS obs, 550 non-AWS obs</description>
<Point>
<coordinates>-89.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -94.5 W</name>
<styleUrl>#ten</styleUrl>
<description>13 AWS obs, 316 non-AWS obs</description>
<Point>
<coordinates>-94.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -95.5 W</name>
<styleUrl>#ten</styleUrl>
<description>6 AWS obs, 116 non-AWS obs</description>
<Point>
<coordinates>-95.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -69.5 W</name>
<styleUrl>#ten</styleUrl>
<description>8 AWS obs, 162 non-AWS obs</description>
<Point>
<coordinates>-69.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -70.5 W</name>
<styleUrl>#ten</styleUrl>
<description>33 AWS obs, 575 non-AWS obs</description>
<Point>
<coordinates>-70.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -71.5 W</name>
<styleUrl>#ten</styleUrl>
<description>31 AWS obs, 576 non-AWS obs</description>
<Point>
<coordinates>-71.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -72.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 386 non-AWS obs</description>
<Point>
<coordinates>-72.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -73.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 247 non-AWS obs</description>
<Point>
<coordinates>-73.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -79.5 W</name>
<styleUrl>#ten</styleUrl>
<description>28 AWS obs, 485 non-AWS obs</description>
<Point>
<coordinates>-79.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -83.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 233 non-AWS obs</description>
<Point>
<coordinates>-83.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -84.5 W</name>
<styleUrl>#ten</styleUrl>
<description>6 AWS obs, 271 non-AWS obs</description>
<Point>
<coordinates>-84.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -90.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 274 non-AWS obs</description>
<Point>
<coordinates>-90.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -93.5 W</name>
<styleUrl>#ten</styleUrl>
<description>14 AWS obs, 330 non-AWS obs</description>
<Point>
<coordinates>-93.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -95.5 W</name>
<styleUrl>#ten</styleUrl>
<description>25 AWS obs, 277 non-AWS obs</description>
<Point>
<coordinates>-95.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -103.5 W</name>
<styleUrl>#ten</styleUrl>
<description>12 AWS obs, 152 non-AWS obs</description>
<Point>
<coordinates>-103.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -113.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 494 non-AWS obs</description>
<Point>
<coordinates>-113.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -114.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 286 non-AWS obs</description>
<Point>
<coordinates>-114.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -116.5 W</name>
<styleUrl>#ten</styleUrl>
<description>79 AWS obs, 2695 non-AWS obs</description>
<Point>
<coordinates>-116.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -71.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 164 non-AWS obs</description>
<Point>
<coordinates>-71.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -72.5 W</name>
<styleUrl>#ten</styleUrl>
<description>15 AWS obs, 456 non-AWS obs</description>
<Point>
<coordinates>-72.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -85.5 W</name>
<styleUrl>#ten</styleUrl>
<description>16 AWS obs, 218 non-AWS obs</description>
<Point>
<coordinates>-85.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -94.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 177 non-AWS obs</description>
<Point>
<coordinates>-94.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -116.5 W</name>
<styleUrl>#ten</styleUrl>
<description>13 AWS obs, 128 non-AWS obs</description>
<Point>
<coordinates>-116.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -121.5 W</name>
<styleUrl>#ten</styleUrl>
<description>16 AWS obs, 281 non-AWS obs</description>
<Point>
<coordinates>-121.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -84.5 W</name>
<styleUrl>#ten</styleUrl>
<description>13 AWS obs, 198 non-AWS obs</description>
<Point>
<coordinates>-84.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -89.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 238 non-AWS obs</description>
<Point>
<coordinates>-89.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>11 AWS obs, 165 non-AWS obs</description>
<Point>
<coordinates>-96.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -110.5 W</name>
<styleUrl>#ten</styleUrl>
<description>5 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-110.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -118.5 W</name>
<styleUrl>#ten</styleUrl>
<description>12 AWS obs, 230 non-AWS obs</description>
<Point>
<coordinates>-118.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -120.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 174 non-AWS obs</description>
<Point>
<coordinates>-120.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -122.5 W</name>
<styleUrl>#ten</styleUrl>
<description>130 AWS obs, 1375 non-AWS obs</description>
<Point>
<coordinates>-122.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -123.5 W</name>
<styleUrl>#ten</styleUrl>
<description>41 AWS obs, 398 non-AWS obs</description>
<Point>
<coordinates>-123.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -92.5 W</name>
<styleUrl>#ten</styleUrl>
<description>39 AWS obs, 387 non-AWS obs</description>
<Point>
<coordinates>-92.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -94.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 247 non-AWS obs</description>
<Point>
<coordinates>-94.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -96.5 W</name>
<styleUrl>#ten</styleUrl>
<description>25 AWS obs, 232 non-AWS obs</description>
<Point>
<coordinates>-96.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>17 AWS obs, 272 non-AWS obs</description>
<Point>
<coordinates>-119.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -124.5 W</name>
<styleUrl>#ten</styleUrl>
<description>9 AWS obs, 93 non-AWS obs</description>
<Point>
<coordinates>-124.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -121.5 W</name>
<styleUrl>#ten</styleUrl>
<description>31 AWS obs, 293 non-AWS obs</description>
<Point>
<coordinates>-121.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -114.5 W</name>
<styleUrl>#ten</styleUrl>
<description>10 AWS obs, 149 non-AWS obs</description>
<Point>
<coordinates>-114.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -116.5 W</name>
<styleUrl>#ten</styleUrl>
<description>7 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-116.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -118.5 W</name>
<styleUrl>#ten</styleUrl>
<description>18 AWS obs, 166 non-AWS obs</description>
<Point>
<coordinates>-118.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -119.5 W</name>
<styleUrl>#ten</styleUrl>
<description>8 AWS obs, 127 non-AWS obs</description>
<Point>
<coordinates>-119.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -123.5 W</name>
<styleUrl>#ten</styleUrl>
<description>44 AWS obs, 541 non-AWS obs</description>
<Point>
<coordinates>-123.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -123.5 W</name>
<styleUrl>#ten</styleUrl>
<description>13 AWS obs, 341 non-AWS obs</description>
<Point>
<coordinates>-123.5,49.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='10-20% AWS'>
<Placemark>
<name>25.5 N, -100.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>8 AWS obs, 53 non-AWS obs</description>
<Point>
<coordinates>-100.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -80.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>56 AWS obs, 433 non-AWS obs</description>
<Point>
<coordinates>-80.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -82.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>91 AWS obs, 602 non-AWS obs</description>
<Point>
<coordinates>-82.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>13 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-95.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -81.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>59 AWS obs, 279 non-AWS obs</description>
<Point>
<coordinates>-81.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>9 AWS obs, 73 non-AWS obs</description>
<Point>
<coordinates>-91.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -82.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>16 AWS obs, 124 non-AWS obs</description>
<Point>
<coordinates>-82.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>75 AWS obs, 398 non-AWS obs</description>
<Point>
<coordinates>-86.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -87.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>142 AWS obs, 668 non-AWS obs</description>
<Point>
<coordinates>-87.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -88.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>33 AWS obs, 253 non-AWS obs</description>
<Point>
<coordinates>-88.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -92.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 113 non-AWS obs</description>
<Point>
<coordinates>-92.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -96.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>67 AWS obs, 366 non-AWS obs</description>
<Point>
<coordinates>-96.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -85.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 98 non-AWS obs</description>
<Point>
<coordinates>-85.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-86.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -89.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>22 AWS obs, 105 non-AWS obs</description>
<Point>
<coordinates>-89.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -104.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>16 AWS obs, 104 non-AWS obs</description>
<Point>
<coordinates>-104.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -109.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>16 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-109.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -88.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>24 AWS obs, 101 non-AWS obs</description>
<Point>
<coordinates>-88.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -90.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 84 non-AWS obs</description>
<Point>
<coordinates>-90.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -92.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-92.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -104.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>13 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-104.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -106.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>56 AWS obs, 322 non-AWS obs</description>
<Point>
<coordinates>-106.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -111.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 175 non-AWS obs</description>
<Point>
<coordinates>-111.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -84.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>103 AWS obs, 596 non-AWS obs</description>
<Point>
<coordinates>-84.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>94 AWS obs, 421 non-AWS obs</description>
<Point>
<coordinates>-86.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -105.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>26 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-105.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -107.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>8 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-107.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -78.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>30 AWS obs, 250 non-AWS obs</description>
<Point>
<coordinates>-78.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -84.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>82 AWS obs, 515 non-AWS obs</description>
<Point>
<coordinates>-84.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -87.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>69 AWS obs, 303 non-AWS obs</description>
<Point>
<coordinates>-87.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -101.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 125 non-AWS obs</description>
<Point>
<coordinates>-101.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -114.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>10 AWS obs, 79 non-AWS obs</description>
<Point>
<coordinates>-114.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -116.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 115 non-AWS obs</description>
<Point>
<coordinates>-116.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -117.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>141 AWS obs, 585 non-AWS obs</description>
<Point>
<coordinates>-117.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -118.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>150 AWS obs, 895 non-AWS obs</description>
<Point>
<coordinates>-118.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -78.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>108 AWS obs, 734 non-AWS obs</description>
<Point>
<coordinates>-78.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -79.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>53 AWS obs, 284 non-AWS obs</description>
<Point>
<coordinates>-79.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -81.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>125 AWS obs, 534 non-AWS obs</description>
<Point>
<coordinates>-81.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -82.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>85 AWS obs, 499 non-AWS obs</description>
<Point>
<coordinates>-82.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -94.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>39 AWS obs, 165 non-AWS obs</description>
<Point>
<coordinates>-94.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -109.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>21 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-109.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -76.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>164 AWS obs, 741 non-AWS obs</description>
<Point>
<coordinates>-76.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -80.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>36 AWS obs, 280 non-AWS obs</description>
<Point>
<coordinates>-80.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>64 AWS obs, 346 non-AWS obs</description>
<Point>
<coordinates>-86.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -88.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>26 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-88.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -90.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 108 non-AWS obs</description>
<Point>
<coordinates>-90.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -96.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>44 AWS obs, 240 non-AWS obs</description>
<Point>
<coordinates>-96.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -100.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-100.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -115.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>60 AWS obs, 311 non-AWS obs</description>
<Point>
<coordinates>-115.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -116.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>43 AWS obs, 274 non-AWS obs</description>
<Point>
<coordinates>-116.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -121.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>113 AWS obs, 524 non-AWS obs</description>
<Point>
<coordinates>-121.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -90.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-90.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 102 non-AWS obs</description>
<Point>
<coordinates>-91.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -93.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 123 non-AWS obs</description>
<Point>
<coordinates>-93.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -104.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>23 AWS obs, 131 non-AWS obs</description>
<Point>
<coordinates>-104.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -120.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>40 AWS obs, 188 non-AWS obs</description>
<Point>
<coordinates>-120.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -82.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 130 non-AWS obs</description>
<Point>
<coordinates>-82.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -85.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>49 AWS obs, 396 non-AWS obs</description>
<Point>
<coordinates>-85.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 122 non-AWS obs</description>
<Point>
<coordinates>-91.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -94.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>69 AWS obs, 463 non-AWS obs</description>
<Point>
<coordinates>-94.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 149 non-AWS obs</description>
<Point>
<coordinates>-95.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -105.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>51 AWS obs, 289 non-AWS obs</description>
<Point>
<coordinates>-105.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -106.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>32 AWS obs, 234 non-AWS obs</description>
<Point>
<coordinates>-106.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -111.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>60 AWS obs, 396 non-AWS obs</description>
<Point>
<coordinates>-111.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -112.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>32 AWS obs, 172 non-AWS obs</description>
<Point>
<coordinates>-112.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -121.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>59 AWS obs, 451 non-AWS obs</description>
<Point>
<coordinates>-121.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -74.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>159 AWS obs, 958 non-AWS obs</description>
<Point>
<coordinates>-74.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -79.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>45 AWS obs, 206 non-AWS obs</description>
<Point>
<coordinates>-79.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -87.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>33 AWS obs, 196 non-AWS obs</description>
<Point>
<coordinates>-87.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -93.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 108 non-AWS obs</description>
<Point>
<coordinates>-93.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>45 AWS obs, 215 non-AWS obs</description>
<Point>
<coordinates>-95.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -101.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>32 AWS obs, 237 non-AWS obs</description>
<Point>
<coordinates>-101.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -103.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>11 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-103.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -119.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>85 AWS obs, 747 non-AWS obs</description>
<Point>
<coordinates>-119.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -72.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>54 AWS obs, 269 non-AWS obs</description>
<Point>
<coordinates>-72.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -85.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>50 AWS obs, 259 non-AWS obs</description>
<Point>
<coordinates>-85.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -87.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>42 AWS obs, 278 non-AWS obs</description>
<Point>
<coordinates>-87.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -114.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 122 non-AWS obs</description>
<Point>
<coordinates>-114.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -115.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 74 non-AWS obs</description>
<Point>
<coordinates>-115.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -117.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>7 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-117.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -77.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>19 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-77.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -78.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>36 AWS obs, 150 non-AWS obs</description>
<Point>
<coordinates>-78.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>58 AWS obs, 414 non-AWS obs</description>
<Point>
<coordinates>-86.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -101.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>12 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-101.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -102.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>12 AWS obs, 78 non-AWS obs</description>
<Point>
<coordinates>-102.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -104.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>36 AWS obs, 179 non-AWS obs</description>
<Point>
<coordinates>-104.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -124.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>13 AWS obs, 86 non-AWS obs</description>
<Point>
<coordinates>-124.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -70.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>95 AWS obs, 655 non-AWS obs</description>
<Point>
<coordinates>-70.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -71.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>457 AWS obs, 1877 non-AWS obs</description>
<Point>
<coordinates>-71.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -72.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>73 AWS obs, 433 non-AWS obs</description>
<Point>
<coordinates>-72.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>22 AWS obs, 154 non-AWS obs</description>
<Point>
<coordinates>-86.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>31 AWS obs, 180 non-AWS obs</description>
<Point>
<coordinates>-91.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -93.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>77 AWS obs, 437 non-AWS obs</description>
<Point>
<coordinates>-93.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -98.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 90 non-AWS obs</description>
<Point>
<coordinates>-98.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -102.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>24 AWS obs, 97 non-AWS obs</description>
<Point>
<coordinates>-102.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -114.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 137 non-AWS obs</description>
<Point>
<coordinates>-114.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -86.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>30 AWS obs, 174 non-AWS obs</description>
<Point>
<coordinates>-86.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -92.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>56 AWS obs, 326 non-AWS obs</description>
<Point>
<coordinates>-92.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -80.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>10 AWS obs, 54 non-AWS obs</description>
<Point>
<coordinates>-80.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -90.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>29 AWS obs, 168 non-AWS obs</description>
<Point>
<coordinates>-90.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -92.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>97 AWS obs, 449 non-AWS obs</description>
<Point>
<coordinates>-92.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>58 AWS obs, 294 non-AWS obs</description>
<Point>
<coordinates>-95.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -104.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>17 AWS obs, 95 non-AWS obs</description>
<Point>
<coordinates>-104.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -106.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>31 AWS obs, 127 non-AWS obs</description>
<Point>
<coordinates>-106.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -123.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>40 AWS obs, 305 non-AWS obs</description>
<Point>
<coordinates>-123.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -87.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 113 non-AWS obs</description>
<Point>
<coordinates>-87.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>26 AWS obs, 110 non-AWS obs</description>
<Point>
<coordinates>-91.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -93.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>121 AWS obs, 545 non-AWS obs</description>
<Point>
<coordinates>-93.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -94.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>68 AWS obs, 348 non-AWS obs</description>
<Point>
<coordinates>-94.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>31 AWS obs, 186 non-AWS obs</description>
<Point>
<coordinates>-95.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -100.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>9 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-100.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -91.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>19 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-91.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -93.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 162 non-AWS obs</description>
<Point>
<coordinates>-93.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -95.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>15 AWS obs, 122 non-AWS obs</description>
<Point>
<coordinates>-95.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -117.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>16 AWS obs, 74 non-AWS obs</description>
<Point>
<coordinates>-117.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -68.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>16 AWS obs, 67 non-AWS obs</description>
<Point>
<coordinates>-68.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -101.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>18 AWS obs, 114 non-AWS obs</description>
<Point>
<coordinates>-101.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -117.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>32 AWS obs, 264 non-AWS obs</description>
<Point>
<coordinates>-117.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -122.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>207 AWS obs, 1667 non-AWS obs</description>
<Point>
<coordinates>-122.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -124.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>15 AWS obs, 110 non-AWS obs</description>
<Point>
<coordinates>-124.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -89.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>27 AWS obs, 116 non-AWS obs</description>
<Point>
<coordinates>-89.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -117.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>22 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-117.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -122.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>92 AWS obs, 801 non-AWS obs</description>
<Point>
<coordinates>-122.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -110.5 W</name>
<styleUrl>#twenty</styleUrl>
<description>3 AWS obs, 21 non-AWS obs</description>
<Point>
<coordinates>-110.5,49.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='20-30% AWS'>
<Placemark>
<name>25.5 N, -77.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>15 AWS obs, 53 non-AWS obs</description>
<Point>
<coordinates>-77.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -82.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>206 AWS obs, 709 non-AWS obs</description>
<Point>
<coordinates>-82.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>27.5 N, -99.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>17 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-99.5,27.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -81.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>270 AWS obs, 1011 non-AWS obs</description>
<Point>
<coordinates>-81.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>68 AWS obs, 218 non-AWS obs</description>
<Point>
<coordinates>-96.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>104 AWS obs, 405 non-AWS obs</description>
<Point>
<coordinates>-97.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -100.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>29 AWS obs, 113 non-AWS obs</description>
<Point>
<coordinates>-100.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>77 AWS obs, 278 non-AWS obs</description>
<Point>
<coordinates>-84.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>103 AWS obs, 315 non-AWS obs</description>
<Point>
<coordinates>-89.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -93.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>69 AWS obs, 264 non-AWS obs</description>
<Point>
<coordinates>-93.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>353 AWS obs, 1406 non-AWS obs</description>
<Point>
<coordinates>-97.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -100.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>15 AWS obs, 57 non-AWS obs</description>
<Point>
<coordinates>-100.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -94.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>68 AWS obs, 216 non-AWS obs</description>
<Point>
<coordinates>-94.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -95.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>24 AWS obs, 85 non-AWS obs</description>
<Point>
<coordinates>-95.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>15 AWS obs, 52 non-AWS obs</description>
<Point>
<coordinates>-96.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>66 AWS obs, 195 non-AWS obs</description>
<Point>
<coordinates>-97.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -111.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>12 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-111.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -85.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>38 AWS obs, 150 non-AWS obs</description>
<Point>
<coordinates>-85.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -94.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>62 AWS obs, 175 non-AWS obs</description>
<Point>
<coordinates>-94.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>199 AWS obs, 769 non-AWS obs</description>
<Point>
<coordinates>-97.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -98.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>40 AWS obs, 118 non-AWS obs</description>
<Point>
<coordinates>-98.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -99.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>33 AWS obs, 107 non-AWS obs</description>
<Point>
<coordinates>-99.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -103.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-103.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -107.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>16 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-107.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -108.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>17 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-108.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -79.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>30 AWS obs, 84 non-AWS obs</description>
<Point>
<coordinates>-79.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -81.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>51 AWS obs, 177 non-AWS obs</description>
<Point>
<coordinates>-81.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -85.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>44 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-85.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -91.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>17 AWS obs, 42 non-AWS obs</description>
<Point>
<coordinates>-91.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -94.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>57 AWS obs, 159 non-AWS obs</description>
<Point>
<coordinates>-94.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -95.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>41 AWS obs, 157 non-AWS obs</description>
<Point>
<coordinates>-95.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>131 AWS obs, 452 non-AWS obs</description>
<Point>
<coordinates>-97.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -80.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>39 AWS obs, 141 non-AWS obs</description>
<Point>
<coordinates>-80.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -86.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>240 AWS obs, 596 non-AWS obs</description>
<Point>
<coordinates>-86.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -88.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>34 AWS obs, 117 non-AWS obs</description>
<Point>
<coordinates>-88.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>59 AWS obs, 181 non-AWS obs</description>
<Point>
<coordinates>-89.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -90.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>9 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-90.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -91.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>26 AWS obs, 94 non-AWS obs</description>
<Point>
<coordinates>-91.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -107.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 58 non-AWS obs</description>
<Point>
<coordinates>-107.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>92 AWS obs, 277 non-AWS obs</description>
<Point>
<coordinates>-84.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -87.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>19 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-87.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>113 AWS obs, 382 non-AWS obs</description>
<Point>
<coordinates>-89.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -93.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>46 AWS obs, 145 non-AWS obs</description>
<Point>
<coordinates>-93.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -105.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>47 AWS obs, 173 non-AWS obs</description>
<Point>
<coordinates>-105.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -108.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>26 AWS obs, 79 non-AWS obs</description>
<Point>
<coordinates>-108.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -75.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>15 AWS obs, 41 non-AWS obs</description>
<Point>
<coordinates>-75.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -77.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>35 AWS obs, 112 non-AWS obs</description>
<Point>
<coordinates>-77.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -79.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>87 AWS obs, 343 non-AWS obs</description>
<Point>
<coordinates>-79.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -81.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>104 AWS obs, 318 non-AWS obs</description>
<Point>
<coordinates>-81.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -83.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>54 AWS obs, 140 non-AWS obs</description>
<Point>
<coordinates>-83.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 45 non-AWS obs</description>
<Point>
<coordinates>-84.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -95.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>164 AWS obs, 498 non-AWS obs</description>
<Point>
<coordinates>-95.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -105.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>39 AWS obs, 130 non-AWS obs</description>
<Point>
<coordinates>-105.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -122.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>8 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-122.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -80.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>57 AWS obs, 145 non-AWS obs</description>
<Point>
<coordinates>-80.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -83.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>43 AWS obs, 122 non-AWS obs</description>
<Point>
<coordinates>-83.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -85.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>24 AWS obs, 63 non-AWS obs</description>
<Point>
<coordinates>-85.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -88.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>64 AWS obs, 192 non-AWS obs</description>
<Point>
<coordinates>-88.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>70 AWS obs, 168 non-AWS obs</description>
<Point>
<coordinates>-89.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -87.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>84 AWS obs, 278 non-AWS obs</description>
<Point>
<coordinates>-87.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>100 AWS obs, 400 non-AWS obs</description>
<Point>
<coordinates>-89.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -90.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>259 AWS obs, 643 non-AWS obs</description>
<Point>
<coordinates>-90.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>28 AWS obs, 68 non-AWS obs</description>
<Point>
<coordinates>-96.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -75.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>358 AWS obs, 1418 non-AWS obs</description>
<Point>
<coordinates>-75.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>365 AWS obs, 927 non-AWS obs</description>
<Point>
<coordinates>-84.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>87 AWS obs, 238 non-AWS obs</description>
<Point>
<coordinates>-89.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -94.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>169 AWS obs, 437 non-AWS obs</description>
<Point>
<coordinates>-94.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -100.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>42 AWS obs, 103 non-AWS obs</description>
<Point>
<coordinates>-100.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -102.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>13 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-102.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -110.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>36 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-110.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -111.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>93 AWS obs, 254 non-AWS obs</description>
<Point>
<coordinates>-111.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -78.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>46 AWS obs, 153 non-AWS obs</description>
<Point>
<coordinates>-78.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -81.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>143 AWS obs, 452 non-AWS obs</description>
<Point>
<coordinates>-81.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -82.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>178 AWS obs, 429 non-AWS obs</description>
<Point>
<coordinates>-82.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -86.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>89 AWS obs, 233 non-AWS obs</description>
<Point>
<coordinates>-86.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>63 AWS obs, 187 non-AWS obs</description>
<Point>
<coordinates>-96.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -102.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 65 non-AWS obs</description>
<Point>
<coordinates>-102.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -109.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>29 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-109.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -110.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-110.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -70.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>124 AWS obs, 472 non-AWS obs</description>
<Point>
<coordinates>-70.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -80.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>117 AWS obs, 314 non-AWS obs</description>
<Point>
<coordinates>-80.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -81.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>335 AWS obs, 820 non-AWS obs</description>
<Point>
<coordinates>-81.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -82.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>136 AWS obs, 326 non-AWS obs</description>
<Point>
<coordinates>-82.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>133 AWS obs, 342 non-AWS obs</description>
<Point>
<coordinates>-84.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -85.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>102 AWS obs, 309 non-AWS obs</description>
<Point>
<coordinates>-85.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -88.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>307 AWS obs, 890 non-AWS obs</description>
<Point>
<coordinates>-88.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>46 AWS obs, 117 non-AWS obs</description>
<Point>
<coordinates>-97.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -100.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 57 non-AWS obs</description>
<Point>
<coordinates>-100.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -109.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>33 AWS obs, 96 non-AWS obs</description>
<Point>
<coordinates>-109.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -110.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>33 AWS obs, 132 non-AWS obs</description>
<Point>
<coordinates>-110.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -76.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>124 AWS obs, 370 non-AWS obs</description>
<Point>
<coordinates>-76.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -82.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>58 AWS obs, 177 non-AWS obs</description>
<Point>
<coordinates>-82.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -83.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>181 AWS obs, 606 non-AWS obs</description>
<Point>
<coordinates>-83.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -84.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>106 AWS obs, 323 non-AWS obs</description>
<Point>
<coordinates>-84.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -85.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>135 AWS obs, 448 non-AWS obs</description>
<Point>
<coordinates>-85.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -90.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>47 AWS obs, 170 non-AWS obs</description>
<Point>
<coordinates>-90.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>32 AWS obs, 97 non-AWS obs</description>
<Point>
<coordinates>-97.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -76.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>101 AWS obs, 280 non-AWS obs</description>
<Point>
<coordinates>-76.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -91.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>78 AWS obs, 237 non-AWS obs</description>
<Point>
<coordinates>-91.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -97.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>8 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-97.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -89.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>86 AWS obs, 271 non-AWS obs</description>
<Point>
<coordinates>-89.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -91.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>34 AWS obs, 109 non-AWS obs</description>
<Point>
<coordinates>-91.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -93.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>252 AWS obs, 749 non-AWS obs</description>
<Point>
<coordinates>-93.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -103.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>84 AWS obs, 282 non-AWS obs</description>
<Point>
<coordinates>-103.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -119.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>14 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-119.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -122.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>49 AWS obs, 173 non-AWS obs</description>
<Point>
<coordinates>-122.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -124.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>34 AWS obs, 111 non-AWS obs</description>
<Point>
<coordinates>-124.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -121.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>70 AWS obs, 189 non-AWS obs</description>
<Point>
<coordinates>-121.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -79.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>11 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-79.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -98.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>15 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-98.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -123.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>59 AWS obs, 178 non-AWS obs</description>
<Point>
<coordinates>-123.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -94.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>45 AWS obs, 178 non-AWS obs</description>
<Point>
<coordinates>-94.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-96.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -116.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>37 AWS obs, 107 non-AWS obs</description>
<Point>
<coordinates>-116.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -103.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>18 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-103.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -96.5 W</name>
<styleUrl>#thirty</styleUrl>
<description>37 AWS obs, 124 non-AWS obs</description>
<Point>
<coordinates>-96.5,50.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='30-40% AWS'>
<Placemark>
<name>26.5 N, -80.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>512 AWS obs, 962 non-AWS obs</description>
<Point>
<coordinates>-80.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -97.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>52 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-97.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>28.5 N, -97.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>75 AWS obs, 131 non-AWS obs</description>
<Point>
<coordinates>-97.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -82.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>126 AWS obs, 219 non-AWS obs</description>
<Point>
<coordinates>-82.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -95.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>472 AWS obs, 887 non-AWS obs</description>
<Point>
<coordinates>-95.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -98.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>312 AWS obs, 509 non-AWS obs</description>
<Point>
<coordinates>-98.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -95.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>234 AWS obs, 496 non-AWS obs</description>
<Point>
<coordinates>-95.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -102.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>36 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-102.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -93.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>18 AWS obs, 29 non-AWS obs</description>
<Point>
<coordinates>-93.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -96.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>327 AWS obs, 726 non-AWS obs</description>
<Point>
<coordinates>-96.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -98.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>36 AWS obs, 77 non-AWS obs</description>
<Point>
<coordinates>-98.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -111.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>186 AWS obs, 366 non-AWS obs</description>
<Point>
<coordinates>-111.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -112.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>220 AWS obs, 483 non-AWS obs</description>
<Point>
<coordinates>-112.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -92.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>73 AWS obs, 151 non-AWS obs</description>
<Point>
<coordinates>-92.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -80.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>216 AWS obs, 451 non-AWS obs</description>
<Point>
<coordinates>-80.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -85.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>154 AWS obs, 286 non-AWS obs</description>
<Point>
<coordinates>-85.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -88.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>108 AWS obs, 165 non-AWS obs</description>
<Point>
<coordinates>-88.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -103.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>12 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-103.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -106.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>325 AWS obs, 662 non-AWS obs</description>
<Point>
<coordinates>-106.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -94.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>230 AWS obs, 479 non-AWS obs</description>
<Point>
<coordinates>-94.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -108.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>32 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-108.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -76.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>150 AWS obs, 330 non-AWS obs</description>
<Point>
<coordinates>-76.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -78.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>94 AWS obs, 161 non-AWS obs</description>
<Point>
<coordinates>-78.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -94.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>148 AWS obs, 300 non-AWS obs</description>
<Point>
<coordinates>-94.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -95.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>118 AWS obs, 197 non-AWS obs</description>
<Point>
<coordinates>-95.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -96.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>55 AWS obs, 99 non-AWS obs</description>
<Point>
<coordinates>-96.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -97.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>268 AWS obs, 540 non-AWS obs</description>
<Point>
<coordinates>-97.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -99.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>26 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-99.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -102.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>35 AWS obs, 78 non-AWS obs</description>
<Point>
<coordinates>-102.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -109.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>36 AWS obs, 74 non-AWS obs</description>
<Point>
<coordinates>-109.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -113.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>84 AWS obs, 163 non-AWS obs</description>
<Point>
<coordinates>-113.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -74.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>13 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-74.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -78.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>250 AWS obs, 392 non-AWS obs</description>
<Point>
<coordinates>-78.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -79.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>33 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-79.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -83.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>31 AWS obs, 62 non-AWS obs</description>
<Point>
<coordinates>-83.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -84.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>115 AWS obs, 235 non-AWS obs</description>
<Point>
<coordinates>-84.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -86.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>81 AWS obs, 149 non-AWS obs</description>
<Point>
<coordinates>-86.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -97.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>135 AWS obs, 226 non-AWS obs</description>
<Point>
<coordinates>-97.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -104.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>231 AWS obs, 521 non-AWS obs</description>
<Point>
<coordinates>-104.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -78.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>151 AWS obs, 334 non-AWS obs</description>
<Point>
<coordinates>-78.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -80.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>39 AWS obs, 91 non-AWS obs</description>
<Point>
<coordinates>-80.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -88.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>54 AWS obs, 116 non-AWS obs</description>
<Point>
<coordinates>-88.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -90.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>32 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-90.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -99.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>75 AWS obs, 114 non-AWS obs</description>
<Point>
<coordinates>-99.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -108.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>45 AWS obs, 79 non-AWS obs</description>
<Point>
<coordinates>-108.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -74.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>1032 AWS obs, 1630 non-AWS obs</description>
<Point>
<coordinates>-74.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -75.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>765 AWS obs, 1320 non-AWS obs</description>
<Point>
<coordinates>-75.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -77.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>148 AWS obs, 223 non-AWS obs</description>
<Point>
<coordinates>-77.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -84.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>164 AWS obs, 350 non-AWS obs</description>
<Point>
<coordinates>-84.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -99.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>44 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-99.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -100.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>41 AWS obs, 64 non-AWS obs</description>
<Point>
<coordinates>-100.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -101.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>30 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-101.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -71.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>361 AWS obs, 674 non-AWS obs</description>
<Point>
<coordinates>-71.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -72.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>599 AWS obs, 1010 non-AWS obs</description>
<Point>
<coordinates>-72.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -74.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>293 AWS obs, 623 non-AWS obs</description>
<Point>
<coordinates>-74.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -83.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>299 AWS obs, 613 non-AWS obs</description>
<Point>
<coordinates>-83.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -92.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>140 AWS obs, 221 non-AWS obs</description>
<Point>
<coordinates>-92.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -74.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>17 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-74.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -75.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>53 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-75.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -77.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>187 AWS obs, 374 non-AWS obs</description>
<Point>
<coordinates>-77.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -85.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>108 AWS obs, 248 non-AWS obs</description>
<Point>
<coordinates>-85.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -88.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>219 AWS obs, 460 non-AWS obs</description>
<Point>
<coordinates>-88.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -89.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>138 AWS obs, 261 non-AWS obs</description>
<Point>
<coordinates>-89.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -75.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>67 AWS obs, 110 non-AWS obs</description>
<Point>
<coordinates>-75.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -88.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>45 AWS obs, 100 non-AWS obs</description>
<Point>
<coordinates>-88.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>45.5 N, -92.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>155 AWS obs, 256 non-AWS obs</description>
<Point>
<coordinates>-92.5,45.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -122.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>128 AWS obs, 227 non-AWS obs</description>
<Point>
<coordinates>-122.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -119.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>40 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-119.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -100.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>18 AWS obs, 33 non-AWS obs</description>
<Point>
<coordinates>-100.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -121.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>17 AWS obs, 33 non-AWS obs</description>
<Point>
<coordinates>-121.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -113.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>38 AWS obs, 58 non-AWS obs</description>
<Point>
<coordinates>-113.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -110.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>27 AWS obs, 51 non-AWS obs</description>
<Point>
<coordinates>-110.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -110.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>16 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-110.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -111.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>30 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-111.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -114.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>107 AWS obs, 197 non-AWS obs</description>
<Point>
<coordinates>-114.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>52.5 N, -101.5 W</name>
<styleUrl>#fourty</styleUrl>
<description>17 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-101.5,52.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='40-50% AWS'>
<Placemark>
<name>25.5 N, -80.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>371 AWS obs, 436 non-AWS obs</description>
<Point>
<coordinates>-80.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -81.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>332 AWS obs, 441 non-AWS obs</description>
<Point>
<coordinates>-81.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -98.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>138 AWS obs, 190 non-AWS obs</description>
<Point>
<coordinates>-98.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -89.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>57 AWS obs, 60 non-AWS obs</description>
<Point>
<coordinates>-89.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -94.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>122 AWS obs, 157 non-AWS obs</description>
<Point>
<coordinates>-94.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -99.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>56 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-99.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -90.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>207 AWS obs, 251 non-AWS obs</description>
<Point>
<coordinates>-90.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -79.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>83 AWS obs, 86 non-AWS obs</description>
<Point>
<coordinates>-79.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -89.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>27 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-89.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -95.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>138 AWS obs, 159 non-AWS obs</description>
<Point>
<coordinates>-95.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -96.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>462 AWS obs, 579 non-AWS obs</description>
<Point>
<coordinates>-96.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>34.5 N, -93.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>50 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-93.5,34.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -90.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>62 AWS obs, 89 non-AWS obs</description>
<Point>
<coordinates>-90.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -114.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>37 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-114.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -104.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>36 AWS obs, 46 non-AWS obs</description>
<Point>
<coordinates>-104.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -114.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>45 AWS obs, 55 non-AWS obs</description>
<Point>
<coordinates>-114.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -75.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>45 AWS obs, 57 non-AWS obs</description>
<Point>
<coordinates>-75.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -79.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>189 AWS obs, 281 non-AWS obs</description>
<Point>
<coordinates>-79.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -84.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>103 AWS obs, 143 non-AWS obs</description>
<Point>
<coordinates>-84.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -101.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>124 AWS obs, 185 non-AWS obs</description>
<Point>
<coordinates>-101.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -103.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 22 non-AWS obs</description>
<Point>
<coordinates>-103.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -114.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>28 AWS obs, 29 non-AWS obs</description>
<Point>
<coordinates>-114.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -76.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>657 AWS obs, 699 non-AWS obs</description>
<Point>
<coordinates>-76.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -98.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>87 AWS obs, 114 non-AWS obs</description>
<Point>
<coordinates>-98.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -99.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>41 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-99.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -100.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>46 AWS obs, 61 non-AWS obs</description>
<Point>
<coordinates>-100.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -113.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-113.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -76.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>1135 AWS obs, 1568 non-AWS obs</description>
<Point>
<coordinates>-76.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -82.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>261 AWS obs, 364 non-AWS obs</description>
<Point>
<coordinates>-82.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -83.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>216 AWS obs, 307 non-AWS obs</description>
<Point>
<coordinates>-83.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -85.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>139 AWS obs, 166 non-AWS obs</description>
<Point>
<coordinates>-85.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -86.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>333 AWS obs, 475 non-AWS obs</description>
<Point>
<coordinates>-86.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -96.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>99 AWS obs, 120 non-AWS obs</description>
<Point>
<coordinates>-96.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -115.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-115.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -73.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>512 AWS obs, 747 non-AWS obs</description>
<Point>
<coordinates>-73.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -76.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>465 AWS obs, 519 non-AWS obs</description>
<Point>
<coordinates>-76.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -83.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>239 AWS obs, 350 non-AWS obs</description>
<Point>
<coordinates>-83.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -73.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>760 AWS obs, 912 non-AWS obs</description>
<Point>
<coordinates>-73.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -76.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>116 AWS obs, 160 non-AWS obs</description>
<Point>
<coordinates>-76.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -87.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>390 AWS obs, 542 non-AWS obs</description>
<Point>
<coordinates>-87.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -78.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>265 AWS obs, 312 non-AWS obs</description>
<Point>
<coordinates>-78.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -87.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>215 AWS obs, 286 non-AWS obs</description>
<Point>
<coordinates>-87.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -88.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>316 AWS obs, 471 non-AWS obs</description>
<Point>
<coordinates>-88.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -87.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>120 AWS obs, 167 non-AWS obs</description>
<Point>
<coordinates>-87.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -87.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>89 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-87.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -88.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>250 AWS obs, 307 non-AWS obs</description>
<Point>
<coordinates>-88.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -121.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 20 non-AWS obs</description>
<Point>
<coordinates>-121.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -120.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>54 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-120.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>47.5 N, -123.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>60 AWS obs, 88 non-AWS obs</description>
<Point>
<coordinates>-123.5,47.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>48.5 N, -124.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-124.5,48.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -95.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>53 AWS obs, 76 non-AWS obs</description>
<Point>
<coordinates>-95.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -100.5 W</name>
<styleUrl>#fifty</styleUrl>
<description>18 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-100.5,51.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='50-60% AWS'>
<Placemark>
<name>25.5 N, -97.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>39 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-97.5,25.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>26.5 N, -82.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>90 AWS obs, 71 non-AWS obs</description>
<Point>
<coordinates>-82.5,26.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -90.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>391 AWS obs, 358 non-AWS obs</description>
<Point>
<coordinates>-90.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -91.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>190 AWS obs, 158 non-AWS obs</description>
<Point>
<coordinates>-91.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -91.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>40 AWS obs, 40 non-AWS obs</description>
<Point>
<coordinates>-91.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -108.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>12 AWS obs, 10 non-AWS obs</description>
<Point>
<coordinates>-108.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>33.5 N, -92.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>35 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-92.5,33.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>35.5 N, -92.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>128 AWS obs, 100 non-AWS obs</description>
<Point>
<coordinates>-92.5,35.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -82.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>270 AWS obs, 200 non-AWS obs</description>
<Point>
<coordinates>-82.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -107.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>28 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-107.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -77.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>493 AWS obs, 412 non-AWS obs</description>
<Point>
<coordinates>-77.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -82.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>43 AWS obs, 31 non-AWS obs</description>
<Point>
<coordinates>-82.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -86.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>35 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-86.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -98.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>90 AWS obs, 72 non-AWS obs</description>
<Point>
<coordinates>-98.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -100.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>163 AWS obs, 138 non-AWS obs</description>
<Point>
<coordinates>-100.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -77.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>1253 AWS obs, 1251 non-AWS obs</description>
<Point>
<coordinates>-77.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -97.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>35 AWS obs, 35 non-AWS obs</description>
<Point>
<coordinates>-97.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -98.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>50 AWS obs, 47 non-AWS obs</description>
<Point>
<coordinates>-98.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -114.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>32 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-114.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -79.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>335 AWS obs, 254 non-AWS obs</description>
<Point>
<coordinates>-79.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -80.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>304 AWS obs, 266 non-AWS obs</description>
<Point>
<coordinates>-80.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -79.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>69 AWS obs, 69 non-AWS obs</description>
<Point>
<coordinates>-79.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -77.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>244 AWS obs, 210 non-AWS obs</description>
<Point>
<coordinates>-77.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -79.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>139 AWS obs, 104 non-AWS obs</description>
<Point>
<coordinates>-79.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>43.5 N, -78.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>148 AWS obs, 148 non-AWS obs</description>
<Point>
<coordinates>-78.5,43.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>44.5 N, -107.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>59 AWS obs, 48 non-AWS obs</description>
<Point>
<coordinates>-107.5,44.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>46.5 N, -82.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>17 AWS obs, 12 non-AWS obs</description>
<Point>
<coordinates>-82.5,46.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -98.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>127 AWS obs, 121 non-AWS obs</description>
<Point>
<coordinates>-98.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -112.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>78 AWS obs, 70 non-AWS obs</description>
<Point>
<coordinates>-112.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -111.5 W</name>
<styleUrl>#sixty</styleUrl>
<description>37 AWS obs, 27 non-AWS obs</description>
<Point>
<coordinates>-111.5,50.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='60-70% AWS'>
<Placemark>
<name>29.5 N, -93.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>37 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-93.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>30.5 N, -94.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>290 AWS obs, 147 non-AWS obs</description>
<Point>
<coordinates>-94.5,30.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>31.5 N, -88.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>19 AWS obs, 11 non-AWS obs</description>
<Point>
<coordinates>-88.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -87.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>182 AWS obs, 119 non-AWS obs</description>
<Point>
<coordinates>-87.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -111.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>11 AWS obs, 5 non-AWS obs</description>
<Point>
<coordinates>-111.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -112.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>57 AWS obs, 37 non-AWS obs</description>
<Point>
<coordinates>-112.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>39.5 N, -77.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>1876 AWS obs, 1128 non-AWS obs</description>
<Point>
<coordinates>-77.5,39.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -75.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>271 AWS obs, 140 non-AWS obs</description>
<Point>
<coordinates>-75.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -98.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>58 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-98.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -112.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>58 AWS obs, 38 non-AWS obs</description>
<Point>
<coordinates>-112.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -113.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>93 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-113.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -97.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>9 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-97.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -112.5 W</name>
<styleUrl>#seventy</styleUrl>
<description>78 AWS obs, 50 non-AWS obs</description>
<Point>
<coordinates>-112.5,51.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='70-80% AWS'>
<Placemark>
<name>31.5 N, -106.5</name>
<styleUrl>#eighty</styleUrl>
<description>217 AWS obs, 66 non-AWS obs</description>
<Point>
<coordinates>-106.5,31.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -96.5</name>
<styleUrl>#eighty</styleUrl>
<description>90 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-96.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -97.5</name>
<styleUrl>#eighty</styleUrl>
<description>313 AWS obs, 129 non-AWS obs</description>
<Point>
<coordinates>-97.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -97.5</name>
<styleUrl>#eighty</styleUrl>
<description>92 AWS obs, 25 non-AWS obs</description>
<Point>
<coordinates>-97.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -100.5</name>
<styleUrl>#eighty</styleUrl>
<description>83 AWS obs, 24 non-AWS obs</description>
<Point>
<coordinates>-100.5,50.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='80-90% AWS'>
<Placemark>
<name>28.5 N, -93.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>18 AWS obs, 4 non-AWS obs</description>
<Point>
<coordinates>-93.5,28.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>29.5 N, -80.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>28 AWS obs, 6 non-AWS obs</description>
<Point>
<coordinates>-80.5,29.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>32.5 N, -87.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>33 AWS obs, 8 non-AWS obs</description>
<Point>
<coordinates>-87.5,32.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -99.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>158 AWS obs, 28 non-AWS obs</description>
<Point>
<coordinates>-99.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -100.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>145 AWS obs, 32 non-AWS obs</description>
<Point>
<coordinates>-100.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -113.5 W</name>
<styleUrl>#ninety</styleUrl>
<description>122 AWS obs, 23 non-AWS obs</description>
<Point>
<coordinates>-113.5,51.5,0</coordinates>
</Point>
</Placemark>
</Folder>
<Folder name='90-100% AWS'>
<Placemark>
<name>24.5 N, -76.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>15 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-76.5,24.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>36.5 N, -110.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>11 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-110.5,36.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>37.5 N, -110.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>11 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-110.5,37.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -117.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>24 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-117.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>38.5 N, -118.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>11 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-118.5,38.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>40.5 N, -116.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>18 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-116.5,40.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>41.5 N, -114.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>14 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-114.5,41.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>42.5 N, -118.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>18 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-118.5,42.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -101.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>7 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-101.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>49.5 N, -111.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>24 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-111.5,49.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -99.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>63 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-99.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>50.5 N, -101.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>57 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-101.5,50.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -99.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>13 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-99.5,51.5,0</coordinates>
</Point>
</Placemark>
<Placemark>
<name>51.5 N, -101.5 W</name>
<styleUrl>#hundred</styleUrl>
<description>45 AWS obs, 0 non-AWS obs</description>
<Point>
<coordinates>-101.5,51.5,0</coordinates>
</Point>
</Placemark>

</Folder>
</Document>
</kml>

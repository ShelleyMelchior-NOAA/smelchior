<markers>
<marker lat=" 71.29" lng="-156.79"
  html='BARROW, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70026.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70026.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 71.32" lng="-156.62"
  html='NORTH SLOPE, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70027.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70027.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 66.89" lng="-162.61"
  html='KOTZEBUE, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70133.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70133.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 66.90" lng="-151.52"
  html='BETTLES, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70174.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70174.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 65.12" lng="-147.48"
  html='CHATANIKA, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70192.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70192.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 66.58" lng="-145.08"
  html='FORT YUKON, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70194.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70194.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 64.51" lng="-165.43"
  html='NOME, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70200.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70200.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 60.79" lng="-161.84"
  html='BETHEL,AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70219.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70219.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 64.73" lng="-156.93"
  html='GALENA, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70222.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70222.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 62.96" lng="-155.60"
  html='MCGRATH, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70231.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70231.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 64.82" lng="-147.88"
  html='FAIRBANKS, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70261.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70261.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 64.00" lng="-145.73"
  html='FORT GREELY, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70267.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70267.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 64.33" lng="-147.65"
  html='BLAIR LAKES RANGE, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70268.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70268.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 61.27" lng="-149.65"
  html='FT RICHARDSON/BRYANT, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70270.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70270.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 61.16" lng="-149.99"
  html='ANCHORAGE, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70273.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70273.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 62.96" lng="-141.94"
  html='NORTHWAY AIRPORT, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70291.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70291.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 63.37" lng="-143.35"
  html='TANACROSS, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70292.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70292.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 57.16" lng="-170.22"
  html='ST. PAUL ISLAND, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70308.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70308.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 55.20" lng="-162.72"
  html='COLD BAY, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70316.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70316.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 58.68" lng="-156.67"
  html='KING SALMON, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70326.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70326.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 57.74" lng="-152.49"
  html='KODIAK, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70350.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70350.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 59.51" lng="-139.67"
  html='YAKUTAT, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70361.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70361.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 55.05" lng="-131.59"
  html='ANNETTE ISLAND, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70398.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70398.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 52.72" lng=" 174.10"
  html='SHEMYA, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70414.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70414.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 51.88" lng="-176.65"
  html='ADAK, AK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_70454.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_70454.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 24.55" lng=" -81.79"
  html='KEY WEST, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72201.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72201.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 25.76" lng=" -80.38"
  html='MIAMI, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72202.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72202.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.48" lng=" -81.70"
  html='JACKSONVILLE, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72206.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72206.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.89" lng=" -80.03"
  html='CHARLESTON, SC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72208.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72208.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.88" lng=" -81.57"
  html='FORT STEWART/WRIGHT, GA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72209.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72209.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 27.71" lng=" -82.40"
  html='TAMPA, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72210.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72210.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.45" lng=" -84.30"
  html='TALLAHASSEE, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72214.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72214.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.36" lng=" -84.57"
  html='ATLANTA, GA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72215.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72215.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.48" lng=" -86.52"
  html='VALPARAISO/EGLIN, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72221.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72221.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.47" lng=" -87.20"
  html='PENSACOLA, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72222.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72222.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.33" lng=" -84.83"
  html='FORT BENNING, GA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72225.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72225.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.18" lng=" -86.78"
  html='BIRMINGHAM, AL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72230.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72230.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.34" lng=" -89.83"
  html='SLIDELL, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72233.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72233.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.32" lng=" -90.08"
  html='JACKSON, MS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72235.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72235.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.10" lng=" -93.20"
  html='FORT POLK, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72239.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72239.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.13" lng=" -93.22"
  html='LAKE CHARLES, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72240.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72240.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.45" lng=" -93.84"
  html='SHREVEPORT, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72248.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72248.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.84" lng=" -97.30"
  html='FORT WORTH, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72249.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72249.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 25.92" lng=" -97.42"
  html='BROWNSVILLE, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72250.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72250.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 27.78" lng=" -97.51"
  html='CORPUS CHRISTI, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72251.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72251.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.10" lng=" -97.33"
  html='FORT HOOD, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72257.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72257.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 29.37" lng="-100.92"
  html='DEL RIO, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72261.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72261.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.94" lng="-102.19"
  html='MIDLAND, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72265.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72265.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.24" lng="-106.22"
  html='WHITE SANDS, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72269.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72269.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.80" lng="-106.40"
  html='EL PASO, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72270.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72270.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.57" lng="-110.33"
  html='FORT HUACHUCA, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72273.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72273.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.23" lng="-110.96"
  html='TUCSON, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72274.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72274.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.45" lng="-111.95"
  html='PHOENIX, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72278.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72278.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.87" lng="-114.33"
  html='YUMA, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72280.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72280.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.82" lng="-115.68"
  html='EL CENTRO NAF, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72281.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72281.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.82" lng="-117.13"
  html='SAN DIEGO/MONTGOMERY, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72290.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72290.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.25" lng="-119.45"
  html='SAN NICOLAS ISLAND, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72291.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72291.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.85" lng="-117.12"
  html='SAN DIEGO, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72293.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72293.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.17" lng=" -79.03"
  html='FAYETTEVILLE/POPE, NC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72303.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72303.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.78" lng=" -76.88"
  html='MOREHEAD CITY, NC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72305.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72305.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.90" lng=" -76.20"
  html='NORFOLK, VA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72308.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72308.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.10" lng=" -79.94"
  html='GREENSBORO, NC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72317.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72317.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.21" lng=" -80.41"
  html='BLACKSBURG, VA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72318.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72318.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.25" lng=" -86.56"
  html='NASHVILLE, TN, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72327.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72327.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.84" lng=" -92.26"
  html='LITTLE ROCK, AR, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72340.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72340.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.65" lng=" -99.27"
  html='ALTUS AFB, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72352.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72352.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.40" lng=" -97.60"
  html='OKLAHOMA CITY/WILL ROGERS, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72353.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72353.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.42" lng=" -97.38"
  html='OKLAHOMA CITY/TINKER, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72354.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72354.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.60" lng=" -98.40"
  html='FORT SILL, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72355.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72355.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.18" lng=" -97.44"
  html='NORMAN, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72357.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72357.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.23" lng="-101.71"
  html='AMARILLO, TX, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72363.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72363.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.87" lng="-106.70"
  html='SANTA TERESA, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72364.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72364.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.04" lng="-106.62"
  html='ALBUQUERQUE, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72365.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72365.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.02" lng="-110.73"
  html='WINSLOW, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72374.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72374.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.23" lng="-111.82"
  html='FLAGSTAFF, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72376.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72376.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.90" lng="-117.92"
  html='EDWARDS AFB, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72381.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72381.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.95" lng="-116.05"
  html='YUCCA FLATS, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72385.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72385.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.05" lng="-115.18"
  html='LAS VEGAS, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72388.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72388.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.12" lng="-119.12"
  html='POINT MUGU NAS, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72391.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72391.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.57" lng="-120.67"
  html='POINT ARGUELLO, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72392.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72392.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.75" lng="-120.57"
  html='VANDENBERG AFB, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72393.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72393.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.90" lng="-120.45"
  html='SANTA MARIA PUBLIC ARPT, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72394.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72394.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.50" lng=" -77.33"
  html='RICHMOND/BYRD, VA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72401.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72401.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.93" lng=" -75.47"
  html='WALLOPS ISLAND, VA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72402.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72402.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.98" lng=" -77.49"
  html='STERLING, VA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72403.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72403.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.28" lng=" -76.40"
  html='PATUXENT RIVER NAS, MD, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72404.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72404.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.03" lng=" -74.32"
  html='LAKEHURST NAS, NJ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72409.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72409.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.90" lng=" -85.97"
  html='FORT KNOX, KY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72424.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72424.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.42" lng=" -83.82"
  html='WILMINGTON, OH, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72426.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72426.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.24" lng=" -93.40"
  html='SPRINGFIELD, MO, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72440.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72440.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.65" lng=" -97.45"
  html='WICHITA, KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72450.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72450.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.76" lng=" -99.97"
  html='DODGE CITY, KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72451.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72451.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.05" lng=" -96.77"
  html='FORT RILEY, KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72455.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72455.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.07" lng=" -95.63"
  html='TOPEKA, KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72456.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72456.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.70" lng="-104.77"
  html='FORT CARSON, CO, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72468.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72468.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.77" lng="-104.87"
  html='DENVER, CO, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72469.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72469.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.12" lng="-108.52"
  html='GRAND JUNCTION, CO, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72476.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72476.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.00" lng="-110.15"
  html='GREEN RIVER, UT, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72477.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72477.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.37" lng="-120.57"
  html='MERCED/CASTLE, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72481.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72481.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.07" lng="-117.08"
  html='TONOPAH, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72485.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72485.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.57" lng="-119.80"
  html='RENO, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72489.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72489.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.74" lng="-122.22"
  html='OAKLAND, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72493.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72493.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.78" lng="-121.85"
  html='CHICO, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72497.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72497.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.87" lng=" -72.86"
  html='UPTON, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72501.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72501.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.25" lng=" -76.92"
  html='WILLIAMSPORT, PA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72514.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72514.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 42.69" lng=" -73.83"
  html='ALBANY, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72518.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72518.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.12" lng=" -76.12"
  html='SYRACUSE, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72519.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72519.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.53" lng=" -80.22"
  html='PITTSBURGH, PA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72520.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72520.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 42.94" lng=" -78.72"
  html='BUFFALO, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72528.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72528.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.98" lng=" -87.90"
  html='CHICAGO/O\'HARE, IL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72530.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72530.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.88" lng=" -91.70"
  html='CEDAR RAPIDS, IA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72545.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72545.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.32" lng=" -96.37"
  html='OMAHA/VALLEY, NE, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72558.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72558.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.13" lng="-100.70"
  html='NORTH PLATTE, NE, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72562.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72562.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.10" lng="-102.98"
  html='SIDNEY, NE, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72563.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72563.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.15" lng="-104.82"
  html='CHEYENNE, WY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72564.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72564.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.77" lng="-111.95"
  html='SALT LAKE CITY, UT, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72572.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72572.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.72" lng="-114.03"
  html='WENDOVER, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72581.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72581.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.86" lng="-115.74"
  html='ELKO, NV, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72582.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72582.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.15" lng="-122.25"
  html='RED BLUFF, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72591.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72591.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 42.38" lng="-122.88"
  html='MEDFORD, OR, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72597.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72597.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 42.70" lng=" -83.47"
  html='WHITE LAKE, MI, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72632.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72632.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.91" lng=" -84.72"
  html='GAYLORD, MI, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72634.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72634.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.50" lng=" -88.11"
  html='GREEN BAY, WI, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72645.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72645.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.85" lng=" -93.56"
  html='CHANHASSEN, MN, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72649.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72649.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.07" lng=" -98.53"
  html='PICKSTOWN, SD, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72652.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72652.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 45.45" lng=" -98.41"
  html='ABERDEEN, SD, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72659.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72659.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.07" lng="-103.21"
  html='RAPID CITY, SD, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72662.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72662.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.07" lng="-108.48"
  html='RIVERTON, WY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72672.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72672.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.57" lng="-116.21"
  html='BOISE, ID, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72681.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72681.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.91" lng="-123.01"
  html='SALEM, OR, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72694.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72694.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 46.87" lng=" -68.01"
  html='CARIBOU, ME, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72712.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72712.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 48.56" lng=" -93.40"
  html='INTERNATIONAL FALLS, MN, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72747.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72747.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 46.77" lng="-100.76"
  html='BISMARCK, ND, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72764.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72764.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 48.21" lng="-106.63"
  html='GLASGOW, MT, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72768.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72768.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 47.46" lng="-111.39"
  html='GREAT FALLS, MT, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72776.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72776.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 47.68" lng="-117.63"
  html='SPOKANE, WA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72786.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72786.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 47.93" lng="-124.56"
  html='QUILLAYUTE, WA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_72797.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_72797.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.60" lng=" -86.62"
  html='REDSTONE ARSENAL, AL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74001.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74001.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.47" lng=" -76.07"
  html='ABERDEEN PROVING GROUNDS, MD, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74002.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74002.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.17" lng="-112.93"
  html='DUGWAY PROVING GROUNDS, UT, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74003.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74003.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.85" lng="-114.40"
  html='YUMA PROVING GROUNDS, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74004.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74004.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.86" lng="-114.03"
  html='YUMA PROVING GROUNDS (TOWER 31, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74005.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74005.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.92" lng="-113.80"
  html='YUMA PROVING GROUNDS (TOWER M), US &lt;br&gt; &lt;a href="./pngs/t120_obs_74006.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74006.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 47.15" lng="-122.48"
  html='TACOMA/MCCHORD, WA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74206.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74206.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 47.08" lng="-122.58"
  html='FORT LEWIS/GRAY, WA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74207.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74207.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 44.05" lng=" -75.73"
  html='FORT DRUM, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74370.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74370.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.89" lng=" -70.26"
  html='GRAY, ME, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74389.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74389.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 43.88" lng=" -69.93"
  html='BRUNSWICK NAS, ME, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74392.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74392.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.61" lng=" -90.58"
  html='DAVENPORT, IA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74455.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74455.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.83" lng=" -85.42"
  html='JEFFERSON PROVING GROUNDS, IN, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74468.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74468.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.78" lng=" -73.77"
  html='NEW YORK/KENNEDY, NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74486.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74486.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 42.47" lng=" -71.28"
  html='HANSCOM FIELD, MA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74490.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74490.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 41.66" lng=" -69.96"
  html='CHATHAM, MA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74494.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74494.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.80" lng=" -73.30"
  html='BROOKHAVEN LAB., NY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74498.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74498.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 37.50" lng="-122.50"
  html='PILAR POINT, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74504.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74504.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.97" lng="-104.82"
  html='U.S. AIR FORCE ACADEMY, CO, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74531.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74531.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.65" lng=" -97.80"
  html='SMOKY HILL GUN. RNG., KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74545.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74545.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 38.62" lng=" -97.30"
  html='HILLSBORO, KS, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74547.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74547.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 40.15" lng=" -89.34"
  html='LINCOLN, IL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74560.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74560.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 39.83" lng=" -84.05"
  html='WRIGHT-PATTERSON AFB, OH, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74570.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74570.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.65" lng="-120.57"
  html='VANDENBERG AFB, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74606.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74606.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.28" lng="-116.62"
  html='BICYCLE LAKE AAF, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74611.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74611.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.68" lng="-117.68"
  html='CHINA LAKE NAF, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74612.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74612.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.27" lng="-117.43"
  html='CUDDLEBACK GUNNERY RANGE, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74618.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74618.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.33" lng="-117.10"
  html='SUPERIOR VALLEY RANGE, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74619.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74619.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.45" lng="-111.95"
  html='PHOENIX, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74626.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74626.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.82" lng="-106.67"
  html='STALLION AAF, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74630.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74630.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.17" lng="-106.48"
  html='W.S.M.R. #32, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74631.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74631.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.30" lng="-103.80"
  html='MELROSE GUNNERY RANGE, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74638.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74638.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.43" lng=" -99.53"
  html='WOODWARD, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74641.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74641.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.61" lng=" -97.49"
  html='LAMONT, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74646.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74646.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.68" lng=" -95.87"
  html='MORRIS, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74650.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74650.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 34.97" lng=" -97.70"
  html='PURCELL, OK, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74651.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74651.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.67" lng=" -87.50"
  html='FORT CAMPBELL, KY, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74671.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74671.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.13" lng=" -78.93"
  html='FORT BRAGG, NC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74693.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74693.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 35.68" lng=" -75.90"
  html='DARE COUNTY RANGE, NC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74695.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74695.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 36.33" lng="-119.93"
  html='LEMOORE NAS, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74702.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74702.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.22" lng="-115.87"
  html='SALTON SEA, CA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74718.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74718.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.93" lng="-112.70"
  html='GILA BEND, AZ, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74724.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74724.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.51" lng="-106.05"
  html='HOLLOMAN AFB, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74732.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74732.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.90" lng="-106.40"
  html='NORTHRUP STRIP, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74733.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74733.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 32.63" lng="-106.40"
  html='W.S.M.R. #39, NM, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74734.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74734.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.32" lng=" -92.55"
  html='ALEXANDRIA/ENGLAND, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74754.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74754.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.18" lng=" -92.63"
  html='CLAIBORNE RANGE, LA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74755.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74755.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.07" lng=" -85.58"
  html='PANAMA CITY/TYNDALL, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74775.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74775.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.42" lng=" -86.68"
  html='HURLBURT AFB, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74777.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74777.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 30.57" lng=" -86.32"
  html='EGLIN AFB RANGE, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74778.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74778.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 31.90" lng=" -81.63"
  html='FORT STEWART, GA, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74780.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74780.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.97" lng=" -80.48"
  html='SHAW AFB, SC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74790.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74790.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 33.85" lng=" -80.48"
  html='POINSETT RANGE, SC, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74792.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74792.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
<marker lat=" 28.47" lng=" -80.55"
  html='CAPE CANAVERAL, FL, US &lt;br&gt; &lt;a href="./pngs/t120_obs_74794.png" target="_blank" &gt;OBS&lt;/a&gt;
     &lt;br&gt; &lt;a href="./pngs/t120_74794.png" target="_blank" &gt;STATS &lt;/a&gt;'
 />
 
</markers>

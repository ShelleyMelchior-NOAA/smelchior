Avg rpts for all dates/cycles: 13481.02
Avg rpts for 00z: 11299.55
Avg rpts for 06z: 16576.55
Avg rpts for 12z: 15692.77
Avg rpts for 18z: 10355.22
Avg AFZA reports for 00z: 998.77
Avg AFZA unique IDs for 00z: 21.88
Avg AFZA0\* reports for 00z: 373.88
Avg AFZA1\* reports for 00z: 0
Avg AFZA2\* reports for 00z: 221.33
Avg AFZA3\* reports for 00z: 0
Avg AFZA4\* reports for 00z: 1.22
Avg AFZA5\* reports for 00z: 15.55
Avg AFZA6\* reports for 00z: 310.55
Avg AFZA7\* reports for 00z: 76.22
Avg AFZA8\* reports for 00z: 0
Avg AFZA9\* reports for 00z: 0
Avg AFZA reports for 06z: 1240.22
Avg AFZA unique IDs for 06z: 34.33
Avg AFZA0\* reports for 06z: 237.88
Avg AFZA1\* reports for 06z: 0
Avg AFZA2\* reports for 06z: 123.88
Avg AFZA3\* reports for 06z: 0
Avg AFZA4\* reports for 06z: 267.55
Avg AFZA5\* reports for 06z: 78.22
Avg AFZA6\* reports for 06z: 217.88
Avg AFZA7\* reports for 06z: 314.77
Avg AFZA8\* reports for 06z: 0
Avg AFZA9\* reports for 06z: 0
Avg AFZA reports for 12z: 1281.00
Avg AFZA unique IDs for 12z: 26.22
Avg AFZA0\* reports for 12z: 190.88
Avg AFZA1\* reports for 12z: 0
Avg AFZA2\* reports for 12z: 71.66
Avg AFZA3\* reports for 12z: 0
Avg AFZA4\* reports for 12z: 394.88
Avg AFZA5\* reports for 12z: 85.88
Avg AFZA6\* reports for 12z: 149.88
Avg AFZA7\* reports for 12z: 387.77
Avg AFZA8\* reports for 12z: 0
Avg AFZA9\* reports for 12z: 0
Avg AFZA reports for 18z: 1156.77
Avg AFZA unique IDs for 18z: 32.11
Avg AFZA0\* reports for 18z: 265.66
Avg AFZA1\* reports for 18z: 0
Avg AFZA2\* reports for 18z: 173.44
Avg AFZA3\* reports for 18z: 0
Avg AFZA4\* reports for 18z: 255.00
Avg AFZA5\* reports for 18z: 40.44
Avg AFZA6\* reports for 18z: 166.11
Avg AFZA7\* reports for 18z: 256.11
Avg AFZA8\* reports for 18z: 0
Avg AFZA9\* reports for 18z: 0
Avg AU reports for 00z: 2727.33
Avg AU unique IDs for 00z: 48.00
Avg AU00\* reports for 00z: 287.33
Avg AU01\* reports for 00z: 2433.66
Avg AU reports for 06z: 2872.33
Avg AU unique IDs for 06z: 49.77
Avg AU00\* reports for 06z: 246.44
Avg AU01\* reports for 06z: 2625.88
Avg AU reports for 12z: 1289.88
Avg AU unique IDs for 12z: 34.22
Avg AU00\* reports for 12z: 252.22
Avg AU01\* reports for 12z: 1037.66
Avg AU reports for 18z: 1065.22
Avg AU unique IDs for 18z: 25.66
Avg AU00\* reports for 18z: 343.11
Avg AU01\* reports for 18z: 702.44
Avg CNC reports for 00z: 184.44
Avg CNC unique IDs for 00z: 2.22
Avg CNCOVM reports for 00z: 107.44
Avg CNCOVL reports for 00z: 21.77
Avg CNCMVT reports for 00z: 55.22
Avg CNCMTS reports for 00z: 0
Avg CNCSVN reports for 00z: 0
Avg CNC reports for 06z: 364.44
Avg CNC unique IDs for 06z: 2.55
Avg CNCOVM reports for 06z: 189.11
Avg CNCOVL reports for 06z: 76.88
Avg CNCMVT reports for 06z: 98.44
Avg CNCMTS reports for 06z: 0
Avg CNCSVN reports for 06z: 0
Avg CNC reports for 12z: 437.55
Avg CNC unique IDs for 12z: 2.88
Avg CNCOVM reports for 12z: 226.88
Avg CNCOVL reports for 12z: 83.66
Avg CNCMVT reports for 12z: 126.77
Avg CNCMTS reports for 12z: .11
Avg CNCSVN reports for 12z: .11
Avg CNC reports for 18z: 129.00
Avg CNC unique IDs for 18z: 2.11
Avg CNCOVM reports for 18z: 68.22
Avg CNCOVL reports for 18z: 18.00
Avg CNCMVT reports for 18z: 42.77
Avg CNCMTS reports for 18z: 0
Avg CNCSVN reports for 18z: 0
Avg CNF reports for 00z: 2327.66
Avg CNF unique IDs for 00z: 27.11
Avg CNFL\* reports for 00z: 511.88
Avg CNFM\* reports for 00z: 0
Avg CNFN\* reports for 00z: 529.77
Avg CNFO\* reports for 00z: 410.11
Avg CNFP\* reports for 00z: 734.00
Avg CNFQ\* reports for 00z: 141.77
Avg CNFR\* reports for 00z: .11
Avg CNF reports for 06z: 4032.88
Avg CNF unique IDs for 06z: 29.33
Avg CNFL\* reports for 06z: 934.88
Avg CNFM\* reports for 06z: .44
Avg CNFN\* reports for 06z: 947.33
Avg CNFO\* reports for 06z: 648.66
Avg CNFP\* reports for 06z: 1289.00
Avg CNFQ\* reports for 06z: 212.55
Avg CNFR\* reports for 06z: 0
Avg CNF reports for 12z: 4038.77
Avg CNF unique IDs for 12z: 29.77
Avg CNFL\* reports for 12z: 932.33
Avg CNFM\* reports for 12z: .33
Avg CNFN\* reports for 12z: 1017.33
Avg CNFO\* reports for 12z: 604.77
Avg CNFP\* reports for 12z: 1232.66
Avg CNFQ\* reports for 12z: 251.11
Avg CNFR\* reports for 12z: .22
Avg CNF reports for 18z: 766.33
Avg CNF unique IDs for 18z: 17.00
Avg CNFL\* reports for 18z: 129.00
Avg CNFM\* reports for 18z: 0
Avg CNFN\* reports for 18z: 229.11
Avg CNFO\* reports for 18z: 91.88
Avg CNFP\* reports for 18z: 262.44
Avg CNFQ\* reports for 18z: 53.88
Avg CNFR\* reports for 18z: 0
Avg EU reports for 00z: 1985.22
Avg EU unique IDs for 00z: 79.88
Avg EU0\* reports for 00z: 1169.77
Avg EU1\* reports for 00z: 185.44
Avg EU2\* reports for 00z: 168.44
Avg EU3\* reports for 00z: 125.44
Avg EU4\* reports for 00z: 55.55
Avg EU5\* reports for 00z: 65.55
Avg EU6\* reports for 00z: 53.00
Avg EU7\* reports for 00z: 54.00
Avg EU8\* reports for 00z: 96.66
Avg EU9\* reports for 00z: 11.33
Avg EU reports for 06z: 4471.11
Avg EU unique IDs for 06z: 155.55
Avg EU0\* reports for 06z: 2601.66
Avg EU1\* reports for 06z: 275.00
Avg EU2\* reports for 06z: 316.66
Avg EU3\* reports for 06z: 269.33
Avg EU4\* reports for 06z: 294.77
Avg EU5\* reports for 06z: 162.22
Avg EU6\* reports for 06z: 164.11
Avg EU7\* reports for 06z: 163.22
Avg EU8\* reports for 06z: 109.22
Avg EU9\* reports for 06z: 114.88
Avg EU reports for 12z: 6803.11
Avg EU unique IDs for 12z: 202.55
Avg EU0\* reports for 12z: 4498.33
Avg EU1\* reports for 12z: 222.77
Avg EU2\* reports for 12z: 355.77
Avg EU3\* reports for 12z: 373.33
Avg EU4\* reports for 12z: 312.33
Avg EU5\* reports for 12z: 189.00
Avg EU6\* reports for 12z: 261.22
Avg EU7\* reports for 12z: 321.88
Avg EU8\* reports for 12z: 86.33
Avg EU9\* reports for 12z: 182.11
Avg EU reports for 18z: 6503.33
Avg EU unique IDs for 18z: 192.44
Avg EU0\* reports for 18z: 4338.55
Avg EU1\* reports for 18z: 265.77
Avg EU2\* reports for 18z: 402.33
Avg EU3\* reports for 18z: 298.44
Avg EU4\* reports for 18z: 319.22
Avg EU5\* reports for 18z: 195.77
Avg EU6\* reports for 18z: 188.66
Avg EU7\* reports for 18z: 226.22
Avg EU8\* reports for 18z: 124.11
Avg EU9\* reports for 18z: 144.22
Avg JP reports for 00z: 2078.88
Avg JP unique IDs for 00z: 171.88
Avg JP9Z4\* reports for 00z: 625.66
Avg JP9Z5\* reports for 00z: 283.44
Avg JP9Z8\* reports for 00z: 62.00
Avg JP9ZV\* reports for 00z: 326.22
Avg JP9ZX\* reports for 00z: 781.55
Avg JP reports for 06z: 2711.55
Avg JP unique IDs for 06z: 196.66
Avg JP9Z4\* reports for 06z: 821.55
Avg JP9Z5\* reports for 06z: 411.55
Avg JP9Z8\* reports for 06z: 77.22
Avg JP9ZV\* reports for 06z: 453.66
Avg JP9ZX\* reports for 06z: 947.55
Avg JP reports for 12z: 1734.77
Avg JP unique IDs for 12z: 180.88
Avg JP9Z4\* reports for 12z: 509.44
Avg JP9Z5\* reports for 12z: 321.88
Avg JP9Z8\* reports for 12z: 38.88
Avg JP9ZV\* reports for 12z: 279.88
Avg JP9ZX\* reports for 12z: 584.66
Avg JP reports for 18z: 153.55
Avg JP unique IDs for 18z: 23.88
Avg JP9Z4\* reports for 18z: 36.33
Avg JP9Z5\* reports for 18z: 63.77
Avg JP9Z8\* reports for 18z: .77
Avg JP9ZV\* reports for 18z: 52.66
Avg JP9ZX\* reports for 18z: 0
Avg NZL reports for 00z: 997.22
Avg NZL unique IDs for 00z: 12.33
Avg NZL00\* reports for 00z: 0
Avg NZL01\* reports for 00z: 145.00
Avg NZL02\* reports for 00z: 255.00
Avg NZL03\* reports for 00z: 2.55
Avg NZL04\* reports for 00z: 181.33
Avg NZL05\* reports for 00z: 413.33
Avg NZL06\* reports for 00z: 0
Avg NZL07\* reports for 00z: 0
Avg NZL08\* reports for 00z: 0
Avg NZL09\* reports for 00z: 0
Avg NZL reports for 06z: 884.00
Avg NZL unique IDs for 06z: 12.11
Avg NZL00\* reports for 06z: 0
Avg NZL01\* reports for 06z: 117.22
Avg NZL02\* reports for 06z: 198.22
Avg NZL03\* reports for 06z: 0
Avg NZL04\* reports for 06z: 175.00
Avg NZL05\* reports for 06z: 393.55
Avg NZL06\* reports for 06z: 0
Avg NZL07\* reports for 06z: 0
Avg NZL08\* reports for 06z: 0
Avg NZL09\* reports for 06z: 0
Avg NZL reports for 12z: 107.33
Avg NZL unique IDs for 12z: 3.66
Avg NZL00\* reports for 12z: 0
Avg NZL01\* reports for 12z: 0
Avg NZL02\* reports for 12z: 88.77
Avg NZL03\* reports for 12z: 0
Avg NZL04\* reports for 12z: 3.77
Avg NZL05\* reports for 12z: 14.77
Avg NZL06\* reports for 12z: 0
Avg NZL07\* reports for 12z: 0
Avg NZL08\* reports for 12z: 0
Avg NZL09\* reports for 12z: 0
Avg NZL reports for 18z: 581.00
Avg NZL unique IDs for 18z: 9.88
Avg NZL00\* reports for 18z: 0
Avg NZL01\* reports for 18z: 92.00
Avg NZL02\* reports for 18z: 125.55
Avg NZL03\* reports for 18z: 0
Avg NZL04\* reports for 18z: 82.33
Avg NZL05\* reports for 18z: 281.11
Avg NZL06\* reports for 18z: 0
Avg NZL07\* reports for 18z: 0
Avg NZL08\* reports for 18z: 0
Avg NZL09\* reports for 18z: 0

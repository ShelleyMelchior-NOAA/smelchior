<!DOCTYPE html PUBLIC "-//w3c//dtd html 4.0 transitional//en">
<html>
<head>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <meta http-equiv="Content-Type" content="text/html; charset=iso-8859-1">


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <meta name="Generator" content="WordPerfect 9">


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <meta name="GENERATOR" content="Mozilla/4.79 [en] (Win98; U) [Netscape]">


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <meta name="Author" content="Dennis Keyser">


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <meta name="Description" content="Last revised 5/30/2001">


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  <title>LIST OF DATA TYPES THAT CAN BE DUMPED</title>
  <meta charset="utf-8">
</head>


<body style="color: rgb(0, 0, 0); background-color: rgb(255, 255, 255);" alink="#ff0000" link="#0000ff" vlink="#551a8b">


















&nbsp;
<br>


















<big>Table 1.a&nbsp;&nbsp; List of valid BUFR data types (last
revised 3/15/2018 <span style="font-style: italic;">-&nbsp;</span></big><big><span style="font-style: italic;">no more updating for
past events expected unless something important later found to be
missed or&nbsp;incorrect</span></big><big><span style="font-style: italic;"></span>).
</big><br>


















<br>


















<br>


















&nbsp; Key for INDICATOR ("IND.") column:<br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-weight: bold;">A - data
type is in BUFR /dcom database and is
available for dumping (in boldface)</span><br>


















&nbsp; &nbsp; &nbsp;<span style="font-style: italic;">A - data type is
temporarily not available for dumping (in italics)</span><br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-style: italic;">F - future
data type, currently not available for dumping (also in italics)<br>


















&nbsp; &nbsp; &nbsp;</span><span style="font-weight: bold;"></span><span style="font-style: italic;"></span><span style="font-style: italic;">O
- data
type obsolete, not available for dumping (also in italics)<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span>P - data type is in /pcom database<span style="font-style: italic;"><br>


















</span>&nbsp;&nbsp;&nbsp;&nbsp; U - data type is in BUFR /dcom database
but currently cannot be dumped<br>


















<br>


















&nbsp; Key for RESTRICTED&nbsp;("RESTR.") column:<br>


















&nbsp;&nbsp;&nbsp;&nbsp; YES - some or all reports&nbsp;in this BUFR
subtype are&nbsp;<a href="http://www.nco.ncep.noaa.gov/sib/restricted_data/restricted_data_pmb/">restricted
with respect&nbsp;to redistribution outside of NCEP for some amount of
time</a><br>


















&nbsp; &nbsp; &nbsp;NO &nbsp;- no data types in this BUFR subtype
are&nbsp;restricted, all are fully available for redistribution outside
of NCEP<br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-style: italic;"></span>&nbsp;&nbsp;&nbsp;
<span style="font-style: italic;"></span><br>


















<p><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <caption><br>


















  </caption><tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="vertical-align: top;" colspan="4">
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      
      <center>BUFR TYPE 0 : SURFACE DATA - LAND</center>


















      </td>


















      <td style="vertical-align: top; text-align: left;">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: top;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">synopr<br>


















      </td>


















      <td style="width: 5%; vertical-align: top; font-family: courier new; font-weight: bold;"><span style="font-size: 10pt;"></span>000<br>


















      </td>


















      <td style="width: 2%; vertical-align: top; font-family: courier new; font-weight: bold;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"></span></span>A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Synoptic
- restricted (WMO Resolution 40) manual and automatic (originating from
WMO SYNOP&nbsp;bulletins) </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>synop<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>001<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><font size="+1"><span style="font-size: 10pt;"></span></font>A<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;">Synoptic
- fixed manual and automatic&nbsp;(originating from WMO
SYNOP&nbsp;bulletins) </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">synopm<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">002<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Synoptic
- mobile manual and automatic (originating from WMO SYNOP
MOBIL&nbsp;bulletins) </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>metar<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>007<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>A<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>Aviation
- METAR<span style="font-size: 10pt;"></span></td>


















      <td style="text-align: left; vertical-align: top;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>prflrs<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>008</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>Surface data from NOAA Profiler
Network (NPN) and Multi-Agency Profiler (MAP) sites<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">shefcm<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">010<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Products
(originally in SHEF format) which are not found in any other
SHEF-format BUFR type/subtype<br>


















      </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;">sheff</td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;">011<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;">A<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;">AFOS
products (precipitation) (originally in SHEF
format) </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>scd<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>012<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>A<br>


















      </td>


















      <td style="font-family: courier new; font-weight: bold; vertical-align: top;"><span style="font-size: 10pt;"></span>Aviation
- supplementary climatological data (SCD)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">nacell</td>


















      <td style="font-family: Courier New; font-style: italic;">020</td>


















      <td style="font-family: Courier New; font-style: italic;">F</td>


















      <td style="font-family: Courier New; font-style: italic;">Wind
energy nacelle, restricted</td>


















      <td style="font-style: italic;">YES</td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">synpbr</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">100</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Synoptic
- restricted (WMO Resolution 40) manual and automatic (originally in
BUFR)</td>


















      <td style="vertical-align: top; text-align: left; font-style: italic;">YES</td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">synopb</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">101</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Synoptic
- fixed manual and automatic&nbsp;(originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">synpmb</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">102</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Synoptic
- mobile manual and automatic (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; font-style: italic;">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-weight: bold; font-style: italic;">


















      <td style="text-align: center; width: 939px; vertical-align: top;" colspan="4">BUFR
TYPE 1 : SURFACE
DATA - SEA</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 939px; vertical-align: top;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; width: 44px; vertical-align: top;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;">ships</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001<br>


















      </td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Ship
- manual and automatic,
restricted (originating from WMO SHIP bulletins)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">dbuoy</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Moored
or drifting buoy (originating in WMO&nbsp;FM-18 format)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">mbuoy</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">003<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Moored
buoy (originating in WMO FM-13 format)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>lcman<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>004<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;"><span style="font-size: 10pt;"></span>CMAN station (originally&nbsp;in CMAN
format)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>tideg<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>005<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;"><span style="font-size: 10pt;"></span>Tide
gauge reports (originally in CREX format) <span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>slpbg<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>006<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-style: italic;"><span style="font-size: 10pt;"></span>Sea
level pressure bogus<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>cstgd<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>007<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span><span style="font-size: 10pt;"></span>A
      </td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-weight: bold;"><span style="font-size: 10pt;"></span>U.S. Coast
Guard reports <span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">tidgcm<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">008<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Tide
gauge reports (originally in CMAN format)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">river<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">009<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">USGS
River/Stream data<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">cmansh</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">010</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">C-MAN
station (originally in SHEF format)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">buoysh</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Buoy
(moored or drifting)&nbsp;(originally in SHEF format) - Note: usually
empty</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">tidgsh</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 939px;">Tide
gauge reports (originally in SHEF format) - Note: usually empty</td>


















      <td style="vertical-align: top; text-align: left; width: 44px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">shipsu</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">013</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-weight: bold;">Ship
- manual and automatic, unrestricted&nbsp;(originating from WMO SHIP
bulletins)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">&lt;tbd&gt;</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">014</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-style: italic;">RVF
river forecast data (originally in SHEF format)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">&lt;tbd&gt;</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">101</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-style: italic;">Ship
- manual and automatic,
restricted (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-style: italic;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">dbuoyb</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">102</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-weight: bold;">Drifting
buoy (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">mbuoyb</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">103</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-weight: bold;">Moored
buoy (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">&lt;tbd&gt;</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">113</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">F</td>


















      <td style="font-family: courier new; vertical-align: top; width: 939px; font-style: italic;">Ship
- manual and automatic, unrestricted&nbsp;(originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 44px; font-style: italic;">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center; width: 936px; vertical-align: top;" colspan="4">BUFR
TYPE 2 :
VERTICAL SOUNDINGS (OTHER THAN SATELLITE)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px;">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 936px; vertical-align: top;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; width: 47px; vertical-align: top;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>raobf<span style="font-size: 10pt;"></span></td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>Rawinsonde
- fixed land (originating from WMO TEMP or PILOT bulletins)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>raobm<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>Rawinsonde
- mobile land&nbsp;(originating from WMO TEMP MOBIL or PILOT MOBIL
bulletins)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>raobs<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>Rawinsonde
- ship&nbsp;(originating from WMO TEMP SHIP or PILOT SHIP bulletins)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>dropw<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">004</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>Dropwinsonde (originating from WMO
TEMP
DROP bulletins)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>pibal<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">005</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>PIBAL&nbsp;(originating from
WMO&nbsp;PILOT,&nbsp;PILOT SHIP or PILOT MOBIL bulletins) <span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">ozonlo<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">006<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">F<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new; width: 936px;">Ozone
soundings, low-resolution (from Met Office)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>prflr<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">007</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-style: italic;"><span style="font-size: 10pt;"></span>NOAA Profiler Network (NPN) winds<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>nxrdw<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">008</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>NEXRAD
Velocity&nbsp;Azimuth Display (VAD) winds decoded from radar coded
message<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>prflrp<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">009</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;"><span style="font-size: 10pt;"></span>Profiler winds originating from PIBALS
(WMO PILOT, PILOT SHIP or PILOT MOBIL bulletins)<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;"><span style="font-size: 10pt;"></span>prflrm<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">010</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-style: italic;"><span style="font-size: 10pt;"></span>NOAA Profiler Network (NPN)&nbsp;spectral moments<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>prflrb<span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;"><span style="font-size: 10pt;"></span>Multi-Agency Profiler (MAP)
and&nbsp;acoustic sounder (SODAR) winds<span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rass<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">RASS
temperatures from <span style="font-weight: normal; font-style: italic;">[NOAA Profiler Network (NPN) - obsolete!]</span> and Multi-Agency
Profilers (MAP)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">prflrj<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-style: italic;">Japanese
Meteorological Agency (JMA) profiler winds<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">prflrh<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">014<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-style: italic;">Other&nbsp;profiler
winds (e.g., from Hong Kong)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">ozonhi<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">015<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new;">F<br>


















      </td>


















      <td style="vertical-align: top; font-style: italic; font-family: courier new; width: 936px;">Ozone
soundings, high-resolution (originally in ASCII format)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-weight: bold;"><span style="font-family: Courier New;">prflre</span><br>


















      </td>


















      <td style="vertical-align: top; font-weight: bold;"><span style="font-family: Courier New;">016</span><br>


















      </td>


















      <td style="vertical-align: top; font-family: Courier New; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: Courier New; width: 936px; font-weight: bold;">European
profiler winds<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-weight: bold;">nxrdw2</td>


















      <td style="vertical-align: top; font-family: Courier New; font-weight: bold;">017</td>


















      <td style="vertical-align: top; font-family: Courier New; font-weight: bold;">A</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-weight: bold;">NEXRAD
Velocity&nbsp;Azimuth Display (VAD)
winds generated from&nbsp;Level II decoder</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-weight: bold; font-family: Times New Roman;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">&lt;tbd&gt;</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">018</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Other
radar Velocity Azimuth Display (VAD) winds (e.g., from Europe, New
Zealand)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">towerr</td>


















      <td style="font-family: Courier New; font-style: italic;">020</td>


















      <td style="font-family: Courier New; font-style: italic;">F</td>


















      <td style="font-family: Courier New; font-style: italic;">Wind
energy tower, restricted</td>


















      <td style="font-style: italic;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">towern</td>


















      <td style="font-family: Courier New; font-style: italic;">021</td>


















      <td style="font-family: Courier New; font-style: italic;">F</td>


















      <td style="font-family: Courier New; font-style: italic;">Wind
energy tower, non-restricted</td>


















      <td style="font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">raobfb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">101</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Rawinsonde
- fixed land (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">raobmb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">102</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Rawinsonde
- mobile land (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">raobsb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">103</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Rawinsonde
- ship (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">dropwb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">104</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Dropwinsonde&nbsp;(originally
in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">pibalb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">105</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">PIBAL&nbsp;(originally
in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">prflpb</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">109</td>


















      <td style="vertical-align: top; font-family: Courier New; font-style: italic;">F</td>


















      <td style="vertical-align: top; width: 936px; font-family: Courier New; font-style: italic;">Profiler
winds originating from PIBALS (originally in BUFR)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-family: Times New Roman; font-style: italic;">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center; width: 936px; vertical-align: top;" colspan="4">BUFR
TYPE 3 :
VERTICAL SOUNDINGS (SATELLITE)</td>


















      <td style="vertical-align: top; text-align: left; width: 47px;">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 936px; vertical-align: top;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; width: 47px; vertical-align: top;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">geost</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-style: italic;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-style: italic;">GOES/NESDIS-processed
5x5 field-of-view soundings/brightness temperatures<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">geosth</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">GOES/NESDIS-processed
1x1 field-of-view cloud data<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">geost1</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">003</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">A</td>


















      <td style="font-family: Courier New; font-weight: bold; width: 936px; vertical-align: top;">GOES/NESDIS-processed
1x1 field-of-view soundings/brightness temperatures</td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">gpsro<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">010<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold; width: 936px;">COSMIC,
CHAMP, GRACE,&nbsp;METOP-2(A)/-1(B)(GRAS),&nbsp;SAC-C,&nbsp;TerraSAR-X
and C/NOFS GPS radio
occultation data<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">tovs</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">101</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">O</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top; width: 936px;">POES/NESDIS-processed
TOVS
soundings/brightness temperatures<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">rtovs</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">102</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">O</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top; width: 936px;">POES/NESDIS-processed
RTOVS
soundings/brightness temperatures<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">atovs</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">104</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">POES/NESDIS-processed
ATOVS
soundings/brightness temperatures<br>


















      </td>


















      <td style="vertical-align: top; text-align: left; width: 47px;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-weight: bold; font-style: italic;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 4 : SINGLE
LEVEL UPPER-AIR DATA (OTHER THAN SATELLITE)</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="width: 10%;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">airep&nbsp;</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Manual
AIREP and Automated Automatic Dependent Surveillance (ADS) aircraft
data (originally in AIREP format) (prior to 10/2009 may have also
included AFWA re-encoded AMDAR and MDCRS reports)</td>


















      <td align="left" valign="top"><span style="font-size: 10pt;"></span><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">pirep</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Manual
PIREP format aircraft data (originally in AIREP format)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">amdar</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
AMDAR&nbsp;aircraft data (originally in AMDAR fromat)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">acars</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">004</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
MDCRS ACARS aircraft
data (from
ARINC) (originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">recco</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">005</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Flight
level reconnaissance aircraft data (originally in RECCO format)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">eadas</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">006</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">European
AMDAR&nbsp;aircraft (E-AMDAR) data (originally
in BUFR)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">acarsa</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">007</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Automated
MDCRS ACARS aircraft data (from ARINC via AFWA) (originally in AIREP
format) <span style="font-size: 10pt;"></span></td>


















      <td style="font-style: italic;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">tamdar<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">008<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Automated
TAMDAR-Mesaba aircraft data (from NOAA/ESRL/GSD MADIS) (originally in
netCDF format)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">camdar<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">009<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
Canadian AMDAR aircraft data (originally in BUFR)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">tmdara</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">010</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A
      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
TAMDAR (all types) aircraft data [from Panasonic (AirDAT)] (originally
in BUFR)</td>


















      <td style="font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">kamdar</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
Korean AMDAR aircraft data (originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">tmdarp</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Automated
TAMDAR-PenAir aircraft data (from NOAA/ESRL/GSD MADIS) (originally in
netCDF format)</td>


















      <td style="font-style: italic;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">tmdarc</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Automated
TAMDAR-Chautauqua&nbsp;aircraft data (from NOAA/ESRL/GSD MADIS)
(originally in netCDF format)</td>


















      <td style="font-style: italic;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">famdar</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">014</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Automated
French&nbsp;AMDAR aircraft data (originally in BUFR)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">hdob</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">015</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">High
Density aircraft observations (HDOB) from reconnaissance aircraft
(originally in HDOBB format)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">amdarb</td>


















      <td style="font-family: Courier New; font-weight: bold;">103</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Automated
AMDAR aircraft data (originally in BUFR)</td>


















      <td style="font-weight: bold;">YES</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 5 : SINGLE
LEVEL UPPER-AIR DATA (SATELLITE)</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-style: italic;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
infrared (long-wave) satellite-derived cloud motion - low density (from
NESDIS
server,
originally in OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
visible satellite-derived cloud motion - low density (from NESDIS
server,
originally in OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
water vapor imager satellite-derived cloud motion - low density (from
NESDIS
server, originally in OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">004</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
picture triplet satellite-derived cloud motion (from NESDIS server,
originally in
OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">005</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
infrared (long-wave) satellite-derived cloud motion - high density
(from NESDIS
server,
originally in OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">006</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
water vapor imager satellite-derived cloud motion (from NESDIS server,
originally
in OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">visuw</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">008</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/UW-CIMSS
visible satellite-derived cloud motion</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">009</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
picture triplet satellite-derived cloud motion (from NESDIS server,
originally in
modified OPARCH format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infus</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">010</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES-15
&amp;&nbsp;down/NESDIS
infrared (long-wave) satellite-derived cloud motion (from NESDIS
server,
originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">h2ius</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES-15
&amp; down/NESDIS
water vapor imager satellite-derived cloud motion (from NESDIS server,
originally
in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">visus</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES-15
&amp; down/NESDIS
visible satellite-derived cloud motion (from NESDIS server, originally
in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ptrus</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
picture triplet satellite-derived cloud motion (from NESDIS server,
originally in
BUFR)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">h2sus</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">014</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES/NESDIS
water vapor sounder satellite-derived cloud motion (from NESDIS server,
originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">015<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O
      <br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
infrared (long-wave) satellite-derived cloud motion (from GTS,
originally in BUFR)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------
      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">016<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
water vapor imager satellite-derived cloud motion (from GTS, originally
in BUFR)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------
      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">017<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
visible satellite-derived cloud motion (from GTS, originally in BUFR)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">018<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GOES/NESDIS
water vapor sounder satellite-derived cloud motion (from GTS,
originally in BUFR)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">3p9us<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">019<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES-15
&amp; down/NESDIS
infrared (short-wave) satellite-derived cloud motion (from NESDIS
server, originally in BUFR)<br>


















      </td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">&lt;tbd&gt;</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">020</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">GOES cloud products above 12,000 feet,&nbsp;supplementary to cloud data in METAR reports (originally in ASCII)</td>




      <td style="font-style: italic; vertical-align: top;">NO</td>




    </tr>




    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">021</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">INSAT/KALPANA/India
infrared (long-wave) satellite-derived cloud motion&nbsp;(originally in
SATOB format)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">022</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">INSAT/KALPANA/India
visible satellite-derived cloud motion&nbsp;(originally in
SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">023</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">INSAT/KALPANA/India
water vapor satellite-derived cloud motion&nbsp;(originally in
SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>




      <td style="font-family: Courier New; font-style: italic;">infin</td>




      <td style="font-family: Courier New; font-style: italic;">024</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">INSAT-3D &amp; up India
infrared (long-wave) satellite-derived cloud motion&nbsp;(originally in BUFR)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>




      <td style="font-family: Courier New; font-style: italic;">visin</td>




      <td style="font-family: Courier New; font-style: italic;">025</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">INSAT-3D &amp; up India
visible satellite-derived cloud motion&nbsp;(originally in BUFR)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>




      <td style="font-family: Courier New; font-style: italic;">h20in</td>




      <td style="font-family: Courier New; font-style: italic;">026</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">INDAT-3D &amp; up India
water vapor satellite-derived cloud motion&nbsp;(originally in BUFR)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">infusr</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">030</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">GOES-16
&amp; up/NESDIS
infrared (long-wave) satellite-derived cloud motion (from NESDIS
server, originally in&nbsp;BUFR)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">h2dusr</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">031</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">GOES-16
&amp; up/NESDIS
water vapor imager deep-layer satellite-derived cloud motion (from
NESDIS server, originally in&nbsp;BUFR)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">visusr</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">032</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">GOES-16
&amp; up/NESDIS
visible satellite-derived cloud motion (from NESDIS server, originally
in BUFR)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">h2tusr</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">034</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">GOES-16
&amp; up/NESDIS
water vapor imager cloud-top satellite-derived cloud motion (from
NESDIS server, originally in&nbsp;BUFR)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">3p9usr</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">039</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">GOES-16
&amp; up/NESDIS
infrared (short-wave) satellite-derived cloud motion (from NESDIS
server, originally in&nbsp;BUFR)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">041</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GMS/MTSAT/JMA
infrared (long-wave) satellite-derived cloud motion - low density
(originally in
SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">042</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GMS/MTSAT/JMA
visible satellite-derived cloud motion - low density (originally in
SATOB format) </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">043</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GMS/MTSAT/JMA
water vapor imager satellite-derived cloud motion - low density
(originally in
SATOB format) </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infja<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">044<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GMS/MTSAT/HIMAWAI/JMA
infrared (long-wave) satellite-derived cloud motion (originally in BUFR)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">visja<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">045<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GMS/MTSAT/HIMAWARI/JMA
visible satellite-derived cloud motion (originally in BUFR)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">h20ja<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">046<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GMS/MTSAT/HIMAWARI/JMA
water vapor imager satellite-derived cloud motion (originally in BUFR) <br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">infjan</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">050</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GMS/NESDIS
infrared (long-wave) satellite-derived cloud motion (originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">h2ijan&nbsp;</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">051</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GMS/NESDIS
water vapor imager satellite-derived cloud motion (originally in BUFR)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">061</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">METEOSAT/EUMETSAT
infrared (long-wave) satellite-derived cloud motion - low density, time
frequency
(originally
in SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">062</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">METEOSAT/EUMETSAT
visible satellite-derived cloud motion - low density, time frequency
(originally
in SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">------<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">063</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">METEOSAT/EUMETSAT
water vapor imager satellite-derived cloud motion - low density, time
frequency
(originally in SATOB format)</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infeu</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">064</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">METEOSAT/EUMETSAT
infrared (long-wave) satellite-derived cloud motion
(originally in BUFR)<span style="font-style: italic;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">viseu</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">065</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">METEOSAT/EUMETSAT
visible satellite-derived cloud motion
(originally in BUFR)<span style="font-style: italic;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">h20eu</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">066</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">METEOSAT/EUMETSAT
water vapor imager satellite-derived cloud motion
(originally in BUFR)<span style="font-style: italic;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infmo<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">070<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">AQUA/TERRA
MODIS infrared (long-wave) satellite-derived cloud motion<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">h20mo<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">071<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">AQUA/<span style="font-weight: normal; font-style: italic;">TERRA</span>
MODIS water vapor imager satellite-derived cloud motion <br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infav</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">080</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NOAA-series/METOP-series
AVHRR infrared (long-wave) satellite-derived cloud motion</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">infvr</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">090</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>
VIIRS&nbsp;infrared (long-wave) satellite-derived cloud motion</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center; width: 936px;" colspan="4">BUFR
TYPE 6 : RADAR
DATA</td>


















      <td style="width: 47px;" align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="width: 10px;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 936px;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle; width: 47px;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">radw30</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind superobs (Level III - NIDS)</td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">radw25<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind superobs (Level II.5 - ORPG)</td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;">rd2w00<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">010<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0000-0059 UTC</td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w01<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0100-0159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w02<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0200-0259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w03<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">013<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0300-0359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w04<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">014<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0400-0459 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w05<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">015<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0500-0559 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w06<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">016<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0600-0659 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w07<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">017<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0700-0759 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w08<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">018<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0800-0859 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w09<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">019<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 0900-0959 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w10<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">020<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1000-1059 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w11<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">021<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1100-1159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w12<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">022<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1200-1259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w13<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">023<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1300-1359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w14<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">024<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1400-1459 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w15<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">025<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1500-1559 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w16<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">026<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1600-1659 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w17<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">027<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1700-1759 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w18<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">028<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1800-1859 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w19<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">029<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 1900-1959 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w20<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">030<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 2000-2059 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w21<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">031<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 2100-2159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w22<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">032<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 2200-2259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2w23<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">033<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
radial wind (Level II - GTS) - 2300-2359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r00<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">040<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0000-0059 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r01<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">041<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0100-0159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r02<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">042<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0200-0259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r03<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">043<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0300-0359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r04<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">044<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0400-0459 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r05<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">045<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0500-0559 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r06<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">046<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0600-0659 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r07<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">047<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0700-0759 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r08<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">048<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0800-0859 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r09<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">049<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 0900-0959 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r10<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">050<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1000-1059 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r11<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">051<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1100-1159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r12<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">052<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1200-1259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r13<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">053<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1300-1359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r14<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">054<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1400-1459 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r15<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">055<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1500-1559 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r16<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">056<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1600-1659 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r17<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">057<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1700-1759 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r18<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">058<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1800-1859 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r19<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">059<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 1900-1959 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-size: 10pt;"></span><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r20<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">060<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 2000-2059 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r21<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">061<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 2100-2159 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r22<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">062<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 2200-2259 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rd2r23<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">063<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold; width: 936px;">NEXRAD
reflectivity (Level II - GTS) - 2300-2359 UTC<br>


















      </td>


















      <td style="width: 47px;" align="left" valign="top"><span style="font-size: 10pt;"></span><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">tldplr</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">070</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">P-3
aircraft Tail Doppler Radar (TDR) radial winds</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr00</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">080</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0000-0059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr01</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">081</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0100-0159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr02</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">082</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0200-0259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr03</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">083</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0300-0359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr04</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">084</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0400-0459 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr05</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">085</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0500-0559 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr06</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">086</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0600-0659 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr07</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">087</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0700-0759 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr08</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">088</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0800-0859 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr09</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">089</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 0900-0959 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr10</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">090</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1000-1059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr11</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">091</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1100-1159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr12</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">092</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1200-1259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr13</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">093</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1300-1359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr14</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">094</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1400-1459 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr15</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">095</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1500-1559 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr16</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">096</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1600-1659 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr17</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">097</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1700-1759 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr18</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">098</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1800-1859 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr19</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">099</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 1900-1959 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr20</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">100</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 2000-2059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr21</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">101</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 2100-2159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr22</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">102</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 2200-2259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcr23</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">103</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar reflectivity - 2300-2359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw00</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">110</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind&nbsp;- 0000-0059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw01</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">111</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0100-0159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw02</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">112</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0200-0259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw03</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">113</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0300-0359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw04</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">114</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0400-0459 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw05</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">115</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0500-0559 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw06</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">116</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0600-0659 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw07</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">117</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0700-0759 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw08</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">118</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0800-0859 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw09</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">119</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 0900-0959 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw10</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">120</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1000-1059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw11</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">121</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1100-1159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw12</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">122</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1200-1259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw13</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">123</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1300-1359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw14</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">124</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1400-1459 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw15</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">125</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1500-1559 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw16</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">126</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1600-1659 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw17</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">127</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1700-1759 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw18</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">128</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1800-1859 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw19</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">129</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 1900-1959 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw20</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">130</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 2000-2059 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw21</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">131</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 2100-2159 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw22</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">132</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 2200-2259 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">rdcw23</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">133</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Canadian
radar radial wind - 2300-2359 UTC</td>


















      <td style="width: 47px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
</span><span style="font-size: 10pt;">
<table style="width: 100%; height: 98px;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center; width: 936px;" colspan="4">BUFR
TYPE 7 :
SYNOPTIC FEATURES</td>


















      <td style="width: 43px;" align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="width: 96px;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 56px;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 25px;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="width: 936px;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle; width: 43px;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; width: 10%;">trpstm</td>


















      <td style="font-family: courier new; vertical-align: top; width: 56px;">000</td>


















      <td style="font-family: courier new; vertical-align: top; width: 25px;">P</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px;">Tropical
storms</td>


















      <td style="width: 43px;" align="left" valign="top"><span style="font-size: 10pt;"></span>NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; width: 10%; font-weight: bold;">ltngsr</td>


















      <td style="font-family: courier new; vertical-align: top; width: 56px; font-weight: bold;">001</td>


















      <td style="font-family: courier new; vertical-align: top; width: 25px; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">National
Lightning Detection Network (NLDN) short-range lightning from Vaisala
via NOAAPORT</td>


















      <td style="width: 43px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; width: 10%; font-weight: bold;">ltnglr</td>


















      <td style="font-family: courier new; vertical-align: top; width: 56px; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; width: 25px; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Long-range
Lightning Dectection Network (LLDN) long-range lightning from Vaisala
via NOAAPORT</td>


















      <td style="width: 43px; font-weight: bold;" align="left" valign="top">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">ltngen</td>


















      <td style="font-family: Courier New; font-weight: bold;">003</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Lightning
data from Earth Networks, Inc. (ENI) Total Lightning Network (ENTLN)</td>


















      <td style="font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; width: 10%; font-weight: bold;">bdyhl2</td>


















      <td style="font-family: courier new; vertical-align: top; width: 56px; font-weight: bold;">021</td>


















      <td style="font-family: courier new; vertical-align: top; width: 25px; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; width: 936px; font-weight: bold;">Boundary
layer height from NEXRAD Level II decoder</td>


















      <td style="width: 43px; font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</span><span style="font-size: 10pt;"><br>


















&nbsp;
<p><a name="1.a.8"></a>
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center; vertical-align: top;" colspan="4">BUFR
TYPE 8 :
PHYSICAL/CHEMICAL CONSTITUENTS</td>


















      <td style="vertical-align: top; text-align: left;">&nbsp;</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td style="vertical-align: top;"><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">osbuv</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-style: italic;">010</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series&nbsp;Solar
Backscatter
UltraViolet
radiances-2 (SBUV-2) nadir profile from NESDIS Version 6 BUFR</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: middle;">osbuv8</td>


















      <td style="font-family: Courier New; font-weight: bold;">011</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">NOAA-series
Solar Backscatter
UltraViolet
radiances-2 (SBUV-2) nadir profile from NESDIS Version 8 BUFR</td>


















      <td style="text-align: left; vertical-align: top;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; text-align: left; font-family: Courier New; font-weight: bold;">gome</td>


















      <td style="vertical-align: top; text-align: left; font-family: Courier New; font-weight: bold;">012</td>


















      <td style="vertical-align: top; text-align: left; font-family: Courier New; font-weight: bold;">A</td>


















      <td style="vertical-align: top; text-align: left; font-family: Courier New; font-weight: bold;">METOP-2(A)/-1(B)&nbsp;Global
Ozone Monitoring Experiment-2
(GOME-2) data </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; text-align: left; font-weight: bold; font-family: Courier New;">omi</td>


















      <td style="vertical-align: top; text-align: left; font-weight: bold; font-family: Courier New;">013</td>


















      <td style="vertical-align: top; text-align: left; font-weight: bold; font-family: Courier New;">A</td>


















      <td style="vertical-align: top; text-align: left; font-weight: bold; font-family: Courier New;">Ozone
Monitoring instrument (OMI)</td>


















      <td style="vertical-align: top; text-align: left; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic; font-weight: bold;"><span style="font-weight: normal;">ompsn6</span></td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">014</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">S-NPP&nbsp;Ozone Mapping and Profiler Suite (OMPS)
nadir profile data (Version 6)</td>


















      <td style="vertical-align: top; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">mls</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">015</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">Microwave
Limb Sounder (MLS) ozone &nbsp;<span style="font-weight: bold; color: rgb(255, 0, 0);">--&gt; temporarily
stopped as of 12z 1/31/2017</span></td>


















      <td style="font-family: Times New Roman; vertical-align: top; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;"><span style="font-style: italic; font-weight: normal;">ompst6</span><br>


















      </td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">016</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold; font-style: italic;">O</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">S-NPP&nbsp;Ozone Mapping and Profiler Suite (OMPS)
total column&nbsp;data (Version 6) plus lat/lon corners&nbsp;</td>


















      <td style="vertical-align: top; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">ompsn8</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">017</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>&nbsp;Ozone Mapping and Profiler Suite (OMPS)
nadir profile data (Version 8)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">ompst8</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">018</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>&nbsp;Ozone Mapping and Profiler Suite (OMPS)
total column&nbsp;data (Version 8)&nbsp;</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-style: italic; vertical-align: top; font-family: courier new;">anowfa<br>


















      </td>


















      <td style="font-style: italic; vertical-align: top; font-family: courier new;">020<br>


















      </td>


















      <td style="font-style: italic; vertical-align: top; font-family: courier new;">O<br>


















      </td>


















      <td style="font-style: italic; vertical-align: top; font-family: courier new;">AIRNOW
ozone data - 1- and 8-hour forward average (delayed)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">anowb1<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">021<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">AIRNOW
ozone data - 1-hour backward average (delayed)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">anowb8<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">022<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">AIRNOW
ozone data - 8-hour backward average (delayed)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">anowrt<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">023<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">AIRNOW
ozone data - 1-hour backward average (realtime - ingested hourly)<br>


















      </td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">anowpm</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">031</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">AIRNOW
particulate data - 1-hour backward average (delayed - ingested daily)</td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">anowp1</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">032</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">A</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">AIRNOW
particulate data - 1-hour backward average (realtime - ingested hourly)</td>


















      <td style="font-weight: bold; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">aodmod</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">041</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">MODIS
Aerosol Optical Depth (AOD) data</td>


















      <td style="vertical-align: top; text-align: left; font-weight: bold;">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















<br>


















&nbsp;
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 12: SURFACE
DATA (SATELLITE)</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;">ssmit</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">DMSP/SSM-I
- processed brightness temperatures</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">ssmip</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">DMSP/SSM-I
- operational products derived at FNMOC (ocean surface wind speed,
total precipitable water, rainfall rate, total cloud water, soil
moisture, ice concentration, ice age, ice edge, skin temperature, snow
depth, rain flag, caluclated surface type)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">gpspw</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">GPS
integrated precipitable water (U.S. only, from GSD)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">gnss</td>


















      <td style="font-family: Courier New; font-weight: bold;">004</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Ground-based
GNSS (GPS, etc.) data (U.S. data from ENI)</td>


















      <td style="font-weight: bold;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ersar</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">005</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ERS/SAR</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-style: italic; font-family: Courier New;">ssmisp</td>


















      <td style="font-style: italic; font-family: Courier New;">006</td>


















      <td style="font-style: italic; font-family: Courier New;">F</td>


















      <td style="font-style: italic; font-family: Courier New;">DMSP/SSM-IS
- operational products derived at FNMOC (ocean surface wind speed,
...)</td>


















      <td style="font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">erswn</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">008</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ERS/scatterometer
winds</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ersal</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">009</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ERS/radar
altimeter data</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">sstnv</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">010</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">O</td>


















      <td style="font-family: courier new; font-style: italic; vertical-align: top;">NAVal
OCEANographic Office (NAVOCEANO)/POES
low-resolution sea surface temperatures</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">sstns</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NESDIS/POES
AVHRR sea surface temperature retrievals,&nbsp;brightness temperatures
and albedo<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">sstnvh</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)/POES
high-resolution AVHRR sea surface temperature
retrievals,&nbsp;brightness
temperatures and albedo</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">trmm</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NASA/Tropical
Rainfall Measuring Mission (TRMM)/TMI) <span style="color: rgb(204, 0, 0);">-- t</span><span style="font-style: italic; color: rgb(204, 0, 0);">he </span><span style="font-style: italic; color: rgb(204, 0, 0);" class="searchword0">TRMM</span><span style="font-style: italic; color: rgb(204, 0, 0);"> satellite ceased
to exist ~&nbsp;4/8/15.</span> </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">sstnvp<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">017<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Physical
retrievals of sea surface temperature generated (by NCEP) from AVHRR
brightness temperatures in BUFR subtype 012 [NAVal
OCEANographic Office (NAVOCEANO)/POES] <br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">sstnsp<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">018<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">Physical
retrievals of sea surface temperature generated (by NCEP) from AVHRR
brightness temperatures in BUFR subtype 011 (NESDIS/POES)<span style="font-size: 10pt;"><br>


















      </span></td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">sstnsg<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">022<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NESDIS/GOES
sea surface temperatures<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">sstvcw</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">023</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">S-NPP/NOAA-20&nbsp;VIIRS sea surface temperatures and radiances - clear sky without land
(NESDIS ACSPO processing) </td>


















      <td style="font-style: italic; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">sstvpw</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">024</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">S-NPP/NOAA-20 VIIRS
sea surface temperatures and radiances - probably clear sky without land (NESDIS
ACSPO processing) </td>


















      <td style="font-style: italic; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">sstvdl</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">025</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">S-NPP/NOAA-20&nbsp;VIIRS
sea surface temperatures and radiances- everything but clear sky and probably
clear sky without land (i.e., others leftover with land)&nbsp;(NESDIS
ACSPO processing) </td>


















      <td style="font-style: italic; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">amsrep<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">031<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">AQUA/AMSR-E
ocean surface products (Level II)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">amsrem</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">034</td>


















      <td style="font-family: Courier New; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: Courier New; font-style: italic;">AQUA/AMSR-E
ocean surface swath products originating from the Multi-Instrument Sea
Surface Temperature (MISST) group at the National Climatic Data Center
(NCDC)</td>


















      <td style="font-family: Times New Roman; vertical-align: top; font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">ssmipn</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">103</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">DMSP/SSM-I
- Neural Net-3 products derived at NCEP (ocean surface wind speed,
total precipitable water, total cloud water, sea-surface temperature)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">ascat</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">122</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">A</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">METOP-2(A)/-1(B)&nbsp;50 KM ASCAT products </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;" align="left" valign="top">&lt;tbd&gt;</td>


















      <td style="font-family: Courier New; font-style: italic;" align="left" valign="top">123</td>


















      <td style="font-family: Courier New; font-style: italic;" align="left" valign="top">F</td>


















      <td style="font-family: Courier New; font-style: italic;" align="left" valign="top">METOP-2(A)/-1(B)&nbsp;25 KM ASCAT products</td>


















      <td style="font-family: Courier New; font-style: italic;" align="left" valign="top"><span style="font-family: Times New Roman;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">qscat</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">137</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">QuikSCAT
products</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">wdsat<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">138<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">WindSat
products from NAVY<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;"><span style="font-size: 10pt;"></span>wdsats</td>


















      <td style="font-family: Courier New; font-style: italic;">139</td>


















      <td style="font-family: Courier New; font-style: italic;">F</td>


















      <td style="font-family: Courier New; font-style: italic;">WindSat
products from NESDIS</td>


















      <td style="font-family: Times New Roman;" align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">lgycld</td>


















      <td style="font-family: Courier New; font-weight: bold;">150</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">GOES/NASA(LANGLEY)-processed
1x1 field-of-view cloud data</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">efclam</td>


















      <td style="font-family: Courier New; font-weight: bold;">160</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">University
of Wisconsin GOES imager effective cloud amount data</td>


















      <td style="font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-style: italic; font-family: Courier New;">&lt;tbd&gt;</td>


















      <td style="font-style: italic; font-family: Courier New;">222</td>


















      <td style="font-style: italic; font-family: Courier New;">F</td>


















      <td style="font-style: italic; font-family: Courier New;">GCOM-W/AMSR2
sea surface temperatures</td>


















      <td style="font-style: italic;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">rscat</td>


















      <td style="font-family: Courier New; font-style: italic;">255</td>


















      <td style="font-family: Courier New; font-style: italic;">O</td>


















      <td style="font-family: Courier New; font-style: italic;"><span style="font-weight: normal;">International Space
Station (ISS) 25 KM RAPIDSCAT
product</span>s&nbsp;<span style="color: rgb(204, 0, 0);">-- instrument died 8/19/2016</span><span style="font-size: 10pt;"><span style="color: rgb(204, 0, 0);"></span><span style="color: rgb(204, 0, 0);" class="searchword0"></span><span style="color: rgb(204, 0, 0);"></span></span></td>


















      <td style="font-style: italic;">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</p>


















</span><span style="font-size: 10pt;">
<p><a name="1.a.21"></a>
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 21 :
RADIANCES (SATELLITE MEASURED)</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-style: italic;">1bhrs2&nbsp;</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-style: italic;">021</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series
(14 and earlier)/HIRS-2
(High resolution
InfraRed Sounder-2)
NCEP-processed brightness temperatures</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">1bmsu</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">022</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series
(14 and earlier)/MSU
(Microwave Sounding
Unit) NCEP-processed brightness temperatures</td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">1bamua</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">023</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NOAA-series
(15 and later)<span style="font-style: italic; color: rgb(0, 0, 0); font-weight: normal;"></span>
and&nbsp;METOP-series /AMSU-A
(Advanced Microwave
Sounding
Unit-A) NCEP-processed brightness temperatures</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">1bamub</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">024</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series
(15-17)<span style="font-weight: normal;"></span>/AMSU-B
(Advanced Microwave
Sounding
Unit-B) NCEP-processed brightness temperatures</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">1bhrs3&nbsp;</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">025</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series
(15-17)<span style="font-weight: normal;"></span>/HIRS-3
(High resolution
InfraRed Sounder-3)
NCEP-processed brightness temperatures</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">1bmhs<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">027<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NOAA-series
(18 and later) and&nbsp;METOP-series /MHS
(Microwave Humidity Sounder) NCEP-processed brightness temperatures<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">1bhrs4<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">028<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NOAA-series
(18 and later) and&nbsp;METOP-series /HIRS-4
(High resolution InfraRed Sounder-4) NCEP-processed brightness
temperatures<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">esamua<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">033<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NOAA-series
(15 and later) and&nbsp;METOP-series /AMSU-A&nbsp;processed brightness
temperatures from&nbsp;Regional ATOVS
Retransmission Services (RARS) [consisting of&nbsp;<em></em>EUMETSAT
ATOVS Retransmis<span style="font-weight: bold;">sion
Service (EARS),&nbsp;Asia-Pacific Regional ATOVS Retransmission&nbsp;
Service&nbsp;(AP-RARS) and&nbsp;South
American Regional ATOVS Retransmission Service (SA-RARS)]</span><br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">esamub<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">034<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA-series
(15-17)/AMSU-B&nbsp;processed brightness temperatures from Regional
ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and South&nbsp;American Regional ATOVS
Retransmission
Service (SA-RARS)]</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">eshrs3<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">035<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-weight: bold;">NOAA-series (15-17)/HIRS-3,
and NOAA-series (18 and later) and METOP_series /HIRS-4&nbsp;processed
brightness temperatures from Regional ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and&nbsp;South
American Regional ATOVS Retransmission Service (SA-RARS)]</span><br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">esmhs</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">036</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">NOAA-series
(18 and later) and METOP-series /MHS&nbsp;processed brightness
temperatures&nbsp;from Regional ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and South American Regional ATOVS
Retransmission Service (SA-RARS)]</td>


















      <td style="vertical-align: top; font-weight: bold; font-family: Times New Roman,Times,serif;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">escris</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">037</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span> Cross-track
Infrared Sounder (CrIS) processed&nbsp;apodized radiances (399
channels)&nbsp;from
Regional ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and South American Regional ATOVS
Retransmission Service (SA-RARS)]</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">esatms</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">038</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>&nbsp;Advanced Technology Microwave Sounder (ATMS)
processed brightness temperatures&nbsp;from Regional ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and South American Regional ATOVS
Retransmission Service (SA-RARS)]</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">esiasi</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">039</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">METOP-series/Infrared
Atmospheric Sounding Interferometer (IASI)
processed radiances from Regional ATOVS
Retransmission Services (RARS) [consisting of EUMETSAT ATOVS
Retransmission&nbsp;Service (EARS), Asia-Pacific Regional ATOVS
Retransmission Service (AP-RARS) and South American Regional ATOVS
Retransmission Service (SA-RARS)] (variable number of channels -
currently 500)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">geoimr</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">041</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">GOES
NESDIS-processed 11x17
field-of-view imager
(clear sky) brightness temperatures<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">sevasr</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">042</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">A</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">METEOSAT Second Generation (MSG)
SEVIRI All
Sky Radiances (ASR) (processed)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">sevcsr</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">043</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">A</td>


















      <td style="font-family: Courier New; font-weight: bold;" align="left" valign="top">METEOSAT Second Generation (MSG)
SEVIRI
Clear Sky Radiances (CSR) (processed)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>




      <td style="font-family: Courier New; font-style: italic;">ahicsr</td>




      <td style="font-family: Courier New; font-style: italic;">044</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">HIMAWARI Clear Sky Radiances (CSR) (processed)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>




      <td style="font-family: Courier New; font-style: italic;">gsrasr</td>




      <td style="font-family: Courier New; font-style: italic;">045</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">GOES-16 &amp; up All Sky Radiances (ASR) (processed)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>




      <td style="font-family: Courier New; font-style: italic;">gsrcsr</td>




      <td style="font-family: Courier New; font-style: italic;">046</td>




      <td style="font-family: Courier New; font-style: italic;">F </td>




      <td style="font-family: Courier New; font-style: italic;">GOES-16 &amp; up Clear Sky Radiances (CSR) (processed)</td>




      <td style="font-style: italic;">NO</td>




    </tr>




    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">avcsam<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">051<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;"><span style="font-style: italic; font-weight: normal;">NOAA-17,</span>
METOP-2(A)/AVHRR
GAC NCEP-processed brightness temperatures - clear and over sea<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">avclam<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">052<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;"><span style="font-style: italic; font-weight: normal;">NOAA-17,</span>
METOP-2(A)/AVHRR
GAC NCEP-processed brightness temperatures - cloud or over land<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">avcspm<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">053<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NOAA-18/AVHRR
GAC NCEP-processed brightness temperatures - clear and over sea<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">avclpm<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">054<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NOAA-18/AVHRR
GAC NCEP-processed brightness temperatures - cloud or over land<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">amuata<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">123<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NOAA-series
(15 and later) and METOP-series /AMSU-A (Advanced Microwave Sounding
Unit-A) NCEP-processed&nbsp;(uncorrected) antenna temperatures<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">ssmisu</td>


















      <td style="font-family: Courier New; font-weight: bold;">201</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">DMSP/SSM-IS
- processed brightness temperatures [Unified Pre-Processor (UPP)]</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">cris</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">202</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP&nbsp;Cross-track
Infrared Sounder (CrIS) apodized radiances (399 channels)</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;"><span style="font-family: Times New Roman;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">atms</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">203</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>&nbsp;Advanced
Technology Microwave Sounder (ATMS)
brightness temperatures</td>


















      <td style="font-family: Times New Roman; vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">viirs</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">204</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">S-NPP/NOAA-20&nbsp;Visible/Infrared
Imager/Radiometer Suite
(VIIRS) radiances</td>


















      <td style="font-style: italic; font-family: Times New Roman; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">crisfs</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">205</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">S-NPP/NOAA-20
Cross-track Infrared Sounder (CrIS) full
spectral radiances (2211 channels)</td>


















      <td style="font-style: italic; vertical-align: top;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">crisf4</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">206</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;"><span style="font-weight: bold;">S-NPP</span>/<span style="font-weight: normal; font-style: italic;">NOAA-20</span>
Cross-track Infrared Sounder (CrIS) full
spectral radiances (431&nbsp;channel subset)</td>


















      <td style="vertical-align: top; font-weight: bold;">NO<br>


















      </td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">crisdb</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">212</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span> Cross-track
Infrared Sounder (CrIS)&nbsp;apodized
radiances (399 channels) - direct broadcast from UW/SSEC</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">atmsdb</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">213</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">S-NPP/<span style="font-weight: normal; font-style: italic;">NOAA-20</span> Advanced
Technology Microwave Sounder (ATMS)
brightness temperatures - direct broadcast from UW/SSEC</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">iasidb
      </td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">239</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">METOP-2(A)/-1(B)&nbsp;Infrared
Atmospheric Sounding Interferometer (IASI) - 1C radiance data (variable
number of channels - currently 616 )- direct broadcast from UW/SSEC</td>


















      <td style="vertical-align: top; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">modair</td>


















      <td style="font-family: Courier New; font-style: italic;">240</td>


















      <td style="font-family: Courier New; font-style: italic;">F</td>


















      <td style="font-family: Courier New; font-style: italic;">MODIS/AIRS
radiance/reflectance data (co-located)</td>


















      <td>NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">mtiasi</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">241</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">A</td>


















      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">METOP-2(A)/-1(B)&nbsp;Infrared
Atmospheric Sounding Interferometer (IASI) - 1C radiance data (variable
number of channels - currently 616)</td>


















      <td style="vertical-align: top; text-align: left;"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">saphir</td>


















      <td style="font-family: Courier New; font-weight: bold;">242</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Megha-Tropiques
SAPHIR L1A2 brightness temperatures</td>


















      <td style="font-weight: bold;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">gmi1cr</td>


















      <td style="font-family: Courier New; font-weight: bold;">246</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">GPM-core/GMI
L1C-R
brightness temperatures</td>


















      <td style="font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">amsr2</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">248</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">GCOM-W/AMSR2
L1B brightness temperatures</td>


















      <td style="font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">airsev</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">249</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; vertical-align: top; font-weight: bold;">AQUA/AIRS,
AMSU-A, HSB processed brightness temperatures - every&nbsp;field-of-view</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">airs<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">250<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">AQUA/AIRS,
AMSU-A, HSB processed brightness temperatures - center field-of-view<br>


















      </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">amsre<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">254<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">AQUA/AMSR-E
processed brightness temperatures<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">airswm<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">255<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">AQUA/AIRS,
AMSU-A, HSB processed brightness temperatures - warmest/clearest
field-of-view<br>


















      </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















<br>


















&nbsp;
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 31 :
OCEANOGRAPHIC DATA</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;">bathy</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">eXpendable BathyThermographs (XBT), thermistor chain moorings [via GTS, originating from WMO&nbsp;FM-63 (BATHY) format]</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">tesac</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">
Conductivity-Temperature-Depth (CTD) probes, Argo profiling floats,
moorings [via GTS, originating from WMO&nbsp;FM-64 (TESAC) format]</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">trkob</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">ThermoSalinoGraphs (TSG)&nbsp;[via GTS, originating from WMO&nbsp;FM-62 (TRACKOB) format]</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">axbt</td>


















      <td style="font-family: Courier New; font-weight: bold;">004</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Airborne
eXpendable BathyThermographs (AXBT) (via GTS,&nbsp;originally in ASCII)</td>


















      <td style="font-family: Times New Roman; font-weight: bold;">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">subpfl</td>


















      <td style="font-family: Courier New; font-weight: bold;">005</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Sub-surface reports from&nbsp;glider profiles, <span style="font-style: italic; font-weight: normal;">Argo profiling&nbsp;floats and other moorings</span>&nbsp;(via GTS, originally in BUFR) </td>


















      <td style="font-weight: bold;">NO</td>


















    </tr>


















    <tr>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">xbtcdt</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">006</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">F</td>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">eXpendable BathyThermographs (XBT), eXpendable Conductivity/Temperature/Depth (XCTD) profiles (originally in BUFR) </td>




      <td style="vertical-align: top;">NO</td>




    </tr>




    <tr>




      <td style="font-family: Courier New; font-style: italic; vertical-align: top;">altkob</td>




      <td style="font-family: Courier New; font-style: italic;">007</td>




      <td style="font-family: Courier New; font-style: italic;">F</td>




      <td style="font-family: Courier New; font-style: italic;">Along-track oceanographic observations&nbsp;(originally in BUFR)</td>




      <td>NO</td>




    </tr>




    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ershal</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA
Laboratory for Satellite Altimetry (NLSA) ERS-2 altimeter Sea Surface
Height Anomaly (SSHA) high-resolution
regional</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">tophal</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA
Laboratory for Satellite Altimetry (NLSA) TOPEX altimeter Sea Surface
Height Anomaly (SSHA) high-resolution
regional</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">toplal</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA
Laboratory for Satellite Altimetry (NLSA) TOPEX altimeter Sea Surface
Height Anomaly (SSHA) low-resolution global</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">gfohal</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">014</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O</td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NOAA
Laboratory for Satellite Altimetry (NLSA) GEOSAT Follow-On (GFO)
altimeter SSHA high-resolution
regional</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">nersal<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">101<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) ERS-2&nbsp;altimeter Sea Surface
Height Anomaly (SSHA)
high-resolution global (via DMZNAS) </td>


















      <td align="left" valign="top"><span style="font-size: 10pt;"></span><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ngfoal<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">102<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) GEOSAT Follow-On (GFO) altimeter Sea
Surface Height Anomaly (SSHA)
high-resolution global (via DMZNAS) </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ntpxal<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">103<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) TOPEX altimeter Sea Surface Height
Anomaly (SSHA) high-resolution
global (via DMZNAS) </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">njsnal<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">104<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) JASON-1 altimeter Sea Surface Height
Anomaly (SSHA)
high-resolution global (via DMZNAS) </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">ngfnal<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">105<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;GEOSAT Follow-On (GFO)
Navy-Interim Geophysical Data Record
(NGDR)&nbsp;altimeter wind/wave (2-day&nbsp;delay) (via DMZNAS) </td>


















      <td align="left" valign="top"><span style="font-style: italic;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">cajsww<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">106<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O
      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">CNES/AVISO
JASON-1 Interim Geophysical Data Record (IGDR)&nbsp;altimeter wind/wave
(2-day delay) (via GTS)<br>


















      </td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">gfofww</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">107</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;GEOSAT Follow-On (GFO) altimeter
wind/wave fast-delivery</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">envsww</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">108</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;ENVISAT
altimeter wind/wave fast delivery (via DMZNAS) <span style="font-size: 10pt;"></span>&nbsp;</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">envsal</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">109</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS)&nbsp;ENVISAT altimeter Sea Surface
Height Anomaly (SSHA)
high-resolution
global (via&nbsp;DMZNAS)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">njsnww</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">110</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;JASON-1 altimeter wind/wave fast
delivery (via&nbsp;DMZNAS)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">------</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">111</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">CNES/AVISO/NESDIS/EUMETSAT
JASON-2 Operational Geophysical Data Record (OGDR)&nbsp;altimeter
wind/wave high-resolution global (1-day
delay) (via server&nbsp;dds.nesdis.noaa.gov)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">njsn2o</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">112</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS)&nbsp;JASON-2 Operational Geophysical
Data Record (OGDR)&nbsp;altimeter Sea Surface Height Anomaly (SSHA)
high-resolution global&nbsp;(1-day delay) (via&nbsp;DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">njsn2i</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">113</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS)&nbsp;JASON-2
Interim Geophysical Data Record (IGDR) altimeter Sea Surface Height
Anomaly (SSHA) high-resolution
global&nbsp;(2-day delay) (via DMZNAS) </td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">njs2ww</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">114</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;JASON-2
altimeter wind/wave fast delivery (via DMZNAS) </td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">cnjsal</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">115</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">CNES/AVISO/NESDIS/EUMETSAT
JASON-2 Operational Geophysical Data Record (OGDR) altimeter Sea
Surface Height Anomaly (SSHA) and&nbsp;wind/wave high-resolution global
(1-day delay) (via GTS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">envavi</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">116</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">O</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">AVISO
SSALTO/DUACS
ENVISAT NRT altimeter Sea Level&nbsp;Anomaly (SLA) high-resolution
global (via server&nbsp;ftp.aviso.oceanobs.com)</td>


















      <td style="font-style: italic;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">ncryal</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">117</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) CRYOSAT-2 altimeter Sea Surface Height Anomaly (SSHA)
high-resolution global&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsarao</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">118</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) Satellite with ARgos and ALtika (SARAL) Operational Geophysical
Data
Record (OGDR) altimeter Sea Surface Height Anomaly (SSHA)
high-resolution global (1-day delay)&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsarai&nbsp;</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">119</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Altimeter Processing System
(ALPS) Satellite with ARgos and ALtika (SARAL) Interim Geophysical Data
Record (IGDR) altimeter Sea Surface Height Anomaly (SSHA)
high-resolution global (2-day delay)&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">ncr2ww</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">120</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;CRYOSAT-2 altimeter wind/wave
fast delivery&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsarww</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">121</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;Satellite with ARgos
and&nbsp;ALtika (SARAL)&nbsp;altimeter wind/wave
fast delivery&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">cnsaal</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">122</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">CNES/AVISO/NESDIS/EUMETSAT
Satellite with ARgos and ALtika (SARAL) Operational Geophysical
Data
Record (OGDR) altimeter Sea Surface Height Anomaly (SSHA)
and wind/wave high-resolution global (1-day delay) (via GTS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">cnc2al</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">123</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">CNES/AVISO/NESDIS/EUMETSAT
CRYOSAT-2&nbsp;Operational Geophysical
Data
Record (OGDR) altimeter Sea Surface Height Anomaly (SSHA)
and wind/wave high-resolution global (1-day delay) (via GTS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">cnj3al</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">124</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">CNES/AVISO/NESDIS/EUMETSAT
JASON-3 Operational Geophysical Data Record (OGDR) altimeter Sea
Surface Height Anomaly (SSHA) and wind/wave high-resolution global
(1-day delay) (via GTS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsjn3o</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">125</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO) Altimeter Processing System
(ALPS)&nbsp;JASON-3 Operational Geophysical Data Record (OGDR)
altimeter Sea Surface Height Anomaly (SSHA) high-resolution global
(1-day delay)&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">njsn3i</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">126</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO) Altimeter Processing System (ALPS)
JASON-3 Interim Geophysical Data Record (IGDR) altimeter Sea Surface
Height Anomaly (SSHA) high-resolution global (2-day delay)&nbsp;(via
DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">njs3ww</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">127</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;JASON-3 altimeter wind/wave fast
delivery&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsn3am</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">128</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;SENTINEL-3A Near Real Time (NRT)
altimeter Sea Surface Height Anomaly (SSHA) high-resolution
global&nbsp;(via
DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsn3as</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">129</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;SENTINEL-3A Slow Time Critical
(STC) altimeter Sea Surface Height Anomaly (SSHA) high-resolution
global&nbsp;(via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">nsn3ww</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">130</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A</td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">NAVal
OCEANographic Office (NAVOCEANO)&nbsp;SENTINEL-3A altimeter
wind/wave&nbsp;fast delivery (via DMZNAS)</td>


















      <td style="font-weight: bold;" align="left" valign="top">NO</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















<br>


















&nbsp;
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr style="font-style: italic; font-weight: bold;">


















      <td style="text-align: center;" colspan="4">BUFR TYPE 255 :
INDICATOR FOR LOCAL USE, WITH SUB-CATEGORY</td>


















      <td align="left" valign="top">&nbsp;</td>


















    </tr>


















    <tr>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">MNEMONIC</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">BUFR</span> <br>


















      <span style="font-size: 9pt;">SUBTYPE</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 9pt;">IND.</span><span style="font-size: 10pt;"></span></td>


















      <td><span style="font-size: 10pt;">DESCRIPTION</span></td>


















      <td style="text-align: left; vertical-align: middle;"><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-size: 10pt;">RESTR.?</span></span></span></td>


















    </tr>


















    <tr>


















      <td style="width: 10%; font-family: courier new; vertical-align: top; font-weight: bold;">msoden</td>


















      <td style="width: 5%; font-family: courier new; vertical-align: top; font-weight: bold;">001</td>


















      <td style="width: 2%; font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO&nbsp;MADIS MESONET feed):&nbsp;Denver Urban Drainage
and Flood Control<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoraw</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">002</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;NFIC Remote
Automatic Weather Stations
(RAWS)</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msowst</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">003</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;MesoWest</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoapr</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">004</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Automatic Position
Reporting
(APR) System Weather Network (citizen weather observers)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msokan</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">005</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Kansas Department of
Transportation</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msofla</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">006</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Florida (FAWN and USF)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoiow</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">007</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Iowa Department of
Transportation</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msomin</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">008</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Minnesota Department
of Transportation</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoawx</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">009</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;"Anything Weather"</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msonos</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">010</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;National Ocean
Service Physical Oceanographic Real-Time System
(NOS-PORTS)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoapg</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">011</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;U.S. Army Aberdeen
Proving
Grounds</td>


















      <td align="left" valign="top"><span style="font-size: 10pt;"></span><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msowfy</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">012</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;"Weather for You"</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">msocob<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">013<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">O<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-style: italic;">Mesonet
data (via NOAA/ESRL/GSD MADIS MESONET feed):&nbsp;NWS COOPerative
Observer program (COOP) <br>


















      </td>


















      <td align="left" valign="top"><span style="font-style: italic;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msohad<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">014<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;NWS
Hydrometeorological Automated Data System (HADS)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoaws<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">015<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;AWS Convergence
Technologies, Inc. (Weather Bug)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoien<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">016<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Iowa Environmental<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msokla<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">017<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Oklahoma Mesonet<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msocol<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">018<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Colorado Department
of Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msowtx<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">019<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;West Texas<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msowis<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">020<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;"><span style="font-size: 10pt;"></span>Mesonet data (via NOAA/NCEP/NCO MADIS
MESONET feed): Wisconsin Department of Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msolju<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">021<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Louisiana State
University and Jackson State University<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">mso470<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">022<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Colorado East
Interstate 470<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msodcn<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">023<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;DC Net (urban
mesonets in Washington, CD and New York City)<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoind<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">024<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Indiana Department of
Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoflt<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">025<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Florida Department of
Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msoalk<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">026<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A<br>


















      </td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed): Alaska Department of
Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">msogeo<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">027<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Georgia Department of
Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">msovir<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">028<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Virginia Department
of Transportation<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">msomca<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">029<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">A<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;Missouri Commercial
Agriculture Weather Network<br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">msothr</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">030</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed):&nbsp;any meso-networks
not in one of the above<br>


















      <small><a href="http://www-sdd.fsl.noaa.gov/MADIS/mesonet_providers.html">click
here</a> to see NOAA/FSL's list of meso-networks</small><br>


















      </td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>










      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">msourb</td>










      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">031</td>










      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">A</td>










      <td style="font-family: Courier New; font-weight: bold; vertical-align: top;">Mesonet
data (via NOAA/NCEP/NCO MADIS URBANET&nbsp; feed): &nbsp;Urbanet (National Mesonet Program Nationwide Network of Networks)</td>










      <td style="font-weight: bold; vertical-align: top;">YES</td>










    </tr>










    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">coopmd</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">101</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Automated
cooperative observer data (via NOAA/NCEP/NCO MADIS COOP feed):&nbsp;New
England Pilot Project (NEPP) and&nbsp;Historical Climatology Network -
Modernization (HCN-M) (replaced "Modernized&nbsp;COOP" - NERON
and Alabama providers, November 2009)<span style="font-size: 10pt;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">coopal</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">102</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">NWS
cooperative observer data (originally in&nbsp;SHEF format): many
different providers, not separated out</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-weight: bold;">msocrn</td>


















      <td style="font-family: Courier New; font-weight: bold;">111</td>


















      <td style="font-family: Courier New; font-weight: bold;">A</td>


















      <td style="font-family: Courier New; font-weight: bold;">Mesonet
data (via NOAA/NCEP/NCO MADIS MESONET feed): Climate Reference Network</td>


















      <td style="font-weight: bold;">YES</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">hydden</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">131</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Hydrological
data (via NOAA/NCEP/NCO MADIS HYDRO feed): Denver Urban Drainage and
Flood Control<span style="font-size: 10pt;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">hydoth</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">160</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Hydrological
data (via NOAA/NCEP/NCO MADIS HYDRO feed):&nbsp;other than Denver Urban
Drainage and Flood Control, not separated out</td>


















      <td align="left" valign="top"><span style="font-weight: bold;">YES</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">snow</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">161</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">A</td>


















      <td style="font-family: courier new; vertical-align: top; font-weight: bold;">Snow
data (via NOAA/NCEP/NCO MADIS snow feed): many different providers, not
separated out <span style="font-size: 10pt;"></span></td>


















      <td align="left" valign="top"><span style="font-weight: bold;">NO</span></td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















<br>


















&nbsp;
</p>


















<hr><br>


















<a name="b"></a><br>


















</span></p>


















<p><br>


















<big>Table 1.b&nbsp;&nbsp; Data group mnemonics used to generate BUFR
dump files in the various NCEP networks.&nbsp; These dump files are
then read by the subsequent PREPBUFR processing steps (last revised
2/5/2018</big><big><span style="font-family: times new roman;"><span style="font-style: italic;"> - not completely up to date!</span>).</span></big><br>


















&nbsp;<br>


















<br>


















<span style="font-family: courier new;">Key for NETWORK ("NET") column
- if&nbsp;</span><span style="font-weight: bold;">BOLDFACE AND
UPPER-CASE</span><span style="font-weight: bold; font-family: courier new;">
</span><span style="font-family: courier new;">indicates the dump file
for this group is read in by the subsequent PREPBUFR processing steps
(although not all of the data may be selected for encoding into
PREPBUFR):</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">A/a - group is dumped in Air Quality
Monitoring (AQM) network</span><br>


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">C/c - group is dumped in CDAS network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">F/f
- group is dumped in GDAS&nbsp;network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">G/g
- group is dumped in GFS&nbsp;network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">H/h
- group is dumped in HOURLY network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; M/m -
group is dumped in RTMA and&nbsp;URMA network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">N/n
- group is dumped in NAM&nbsp;network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-style: italic; font-family: courier new;">o &nbsp; - group
is
obsolete and is not dumped in any network (also in italics)</span><br>


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; R/r -
group is dumped in&nbsp;RAP network</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;"></span><span style="font-family: courier new;"></span><span style="font-family: courier new;"></span><span style="font-style: italic; font-family: courier new;"></span><span style="font-family: courier new;"></span><span style="font-style: italic; font-family: courier new;">t &nbsp; - group
consists of future data types and is currently not dumped in any
network (also in italics)</span><br style="font-family: courier new;">


















</p>


















<p><br style="font-family: courier new;">


















<span style="font-family: courier new;">Key for superscripts in "NET"
column:<a name="b.2"></a></span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 1 -
input to QuikSCAT reprocessing program WAVE_DCODQUIKSCAT which outputs
superobed data (on a 0.5 degree lat/lon grid) in a file called
&ldquo;qkswnd&rdquo;
which is read by the subsequent PREPBUFR processing steps if network is
</span><span style="font-weight: bold; font-family: courier new;">boldface<a name="b.1"></a></span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 2 -
input to SSM/I reprocessing program PREPOBS_PREPSSMI which outputs
superobed data (on a 1 degree lat/lon grid) in a file called "spssmi"
which is read by the subsequent PREPBUFR processing steps if network is
</span><span style="font-weight: bold; font-family: courier new;">boldface
</span><span style="font-family: courier new;">[in the GFS and GDAS
networks, the superobed FNMOC rainfall rate product in
&ldquo;spssmi&rdquo; is
currently also read by the Global GSI analysis (the analysis does not
read these data from the PREPBUFR file even though they are written
there)]</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 3 -
input to SSM/I reprocessing program PREPOBS_PREPSSMI which outputs
non-superobed data in a file called "spssmi" which is read by the
subsequent PREPBUFR processing steps if network is </span><span style="font-weight: bold; font-family: courier new;">boldface<br>


















&nbsp;&nbsp;&nbsp;&nbsp; </span><span style="font-family: courier new;">4
- <span style="font-style: italic;">(reserved for future use)</span> </span><span style="font-weight: bold; font-family: courier new;"><a name="b.3"></a></span><br>


















<span style="font-family: courier new;">
&nbsp; &nbsp; &nbsp;5 -&nbsp;</span><span style="font-family: courier new;">input to WindSat&nbsp;reprocessing
program BUFR_DCODWINDSAT which outputs
superobed data (on a 1 degree lat/lon grid) in a file called
&ldquo;wdsatr&rdquo;
which is read by the subsequent PREPBUFR processing steps if network is
</span><span style="font-weight: bold; font-family: courier new;">boldface</span><br>


















<span style="font-family: courier new;">&nbsp; &nbsp; &nbsp;6 -&nbsp;</span><span style="font-family: courier new;">input to WindSat&nbsp;reprocessing
program BUFR_DCODWINDSAT which outputs&nbsp;data (not superobed) in a
file called
&ldquo;wdsatr&rdquo;
which is read by the subsequent PREPBUFR processing steps if network is
</span><span style="font-weight: bold; font-family: courier new;">boldface</span><br>


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 7 -
input to ASCAT&nbsp;reprocessing program WAVE_DCODQUIKSCAT which
outputs&nbsp;data (not superobed) in a file called &ldquo;ascatw&rdquo;
which is read by the subsequent PREPBUFR processing steps if network is
</span><span style="font-weight: bold; font-family: courier new;">boldface<a name="b.6"></a></span><br>


















<span style="font-family: courier new;">&nbsp; &nbsp; &nbsp;8 - even
though this dump file is read&nbsp;by the PREPBUFR processing steps in
this network, the subsequent&nbsp;analysis code reads the same dump
file directly (ignoring&nbsp;the data encoded&nbsp;in the PREPBUFR file
from this dump file)</span></p>


















<p><span style="font-family: courier new;"> </span><br>


















<span style="font-family: courier new;">Key for superscripts in
"MNEMONICS INCLUDED" column:</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 1 -
not included in&nbsp;RAP network dumps</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 2 -
not included in CDAS network dumps</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 3 -
not included in NAM&nbsp;network dumps</span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 4 -
<span style="font-style: italic;">(reserved for future use)</span></span><br style="font-family: courier new;">


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; 5 -
not included in GFS or GDAS network dumps<br>


















&nbsp; &nbsp;&nbsp; 6 - not included in HOURLY network dumps<br>


















&nbsp; &nbsp; &nbsp;7 - included in NAM&nbsp;network dumps but not
read by subsequent PREPBUFR processing steps in these networks <br>


















&nbsp; &nbsp; &nbsp;8 - included in CDAS&nbsp;network dump but
not&nbsp;read by subsequent PREPBUFR processing steps </span><span style="font-family: courier new;">in this network</span><br>


















<span style="font-family: courier new;">
&nbsp; &nbsp; &nbsp;9 - if "acars" contains more reports than "acarsa"
(normally the case) then only "acars" is read by subsequent PREPBUFR
processing steps in all indicated networks<br>


















&nbsp; &nbsp; 10 - </span><span style="font-family: courier new;">if
"acarsa" contains more
reports than "acars" (normally not the case) then only "acarsa" is read
by
subsequent PREPBUFR processing steps in all indicated networks<br>


















&nbsp;&nbsp;&nbsp; 11 -
not included in RTMA and&nbsp;URMA network dumps<br>


















&nbsp; &nbsp; 12 - Not read by subsequent PREPBUFR processing steps in
any network<br>


















&nbsp; &nbsp;&nbsp;13 - Currently only reports from ENI (mainly over
U.S.) are encoded into PREPBUFR file (for every network).&nbsp;
European GNSS reports are skipped.</span><span style="font-size: 10pt;">
<p><br>


















&nbsp;
<table border="1" width="100%">


















  <tbody>


















    <tr valign="top">


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 10pt;"></span><span style="font-size: 10pt;">GROUP
MNEMONIC</span> <br>


















      <span style="font-size: 10pt;">(dump file)</span></td>


















      <td><span style="font-size: 10pt;">NET</span></td>


















      <td><span style="font-size: 10pt;">MNEMONICS INCLUDED (<span style="text-decoration: underline;">underlined</span> means some or
all reports in this mnemonic&nbsp;are <a href="http://www.nco.ncep.noaa.gov/sib/restricted_data/restricted_data_pmb/">restricted
with respect to redistribution outside of NCEP for some amount of time</a>)</span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">adpsfc</span><span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">C</span>,<span style="font-weight: bold;">M</span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;"><span style="font-family: courier new; text-decoration: underline;">synopr</span>,
synop</span><span style="font-family: Courier New;">,
synopm<sup>1,3,11</sup>, metar</span><span style="font-family: Courier New;"></span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">adpupa</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: courier new;"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">C</span></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">raobf,
raobm, raobs, dropw, pibal, recco</span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">aircar</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-weight: bold; font-family: courier new;">R</span><span style="font-family: courier new;">,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">C</span></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;"><span style="text-decoration: underline;">acars</span><sup>9,10</sup>, <span style="text-decoration: underline;">acarsa</span><sup>9,10</sup></span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">aircft</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: courier new;"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">C</span></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">airep,
pirep, <span style="text-decoration: underline;">asdar</span>, <span style="text-decoration: underline;">eadas</span>, <span style="text-decoration: underline;">camdar</span><sup>8</sup> <span style="text-decoration: underline;"></span><span style="text-decoration: underline;"></span><span style="text-decoration: underline;"></span><span style="text-decoration: underline;">tmdara</span><sup>8</sup>,&nbsp;<span style="text-decoration: underline;"></span><span style="text-decoration: underline;">kamdar</span>, <span style="text-decoration: underline;">amdarb</span></span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">airnow<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">A</span><br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">anowb1,
anowb8<br>


















      </td>


















    </tr>


















    <tr valign="top">


















      <td style="font-family: courier new; color: rgb(0, 0, 0);">atovs</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);">f,<span style="font-weight: bold;">C</span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);">atovs</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;" align="left" valign="top">ascatt</td>


















      <td style="font-family: Courier New;" align="left" valign="top"><span style="font-weight: bold;">R<sup>7</sup></span>,<span style="font-weight: bold;">N<sup>7</sup></span>,<span style="font-weight: bold;">G</span><sup style="font-weight: bold;">7</sup>,<span style="font-weight: bold;">F</span><sup style="font-weight: bold;">7</sup>,c<sup>7</sup>,<span style="font-weight: bold;">M</span><sup style="font-weight: bold;">7</sup></td>


















      <td style="font-family: Courier New;" align="left" valign="top">ascat</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">erswnd</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">o<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">erswn</td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">goesnd</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: courier new;"><span style="font-weight: bold;">R,n</span><span style="font-weight: bold;"></span></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">geost1</span><sup><span style="font-size: 10pt;"><span style="font-family: Courier New;">3</span></span></sup><span style="font-family: Courier New;">,
geosth</span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">gpsipw</td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R,N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">gnss<span style="font-size: 10pt;"><sup><span style="font-size: 10pt;"><span style="font-family: Courier New;">13</span></span></sup><span style="font-family: Courier New;"></span></span></td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">msonet</td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R,N</span>,c,<span style="font-weight: bold;">M</span></td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="text-decoration: underline;">msoden</span>, <span style="text-decoration: underline;">msoraw</span>, <span style="text-decoration: underline;">msowst</span>, <span style="text-decoration: underline;">msoapr</span>, <span style="text-decoration: underline;">msokan</span>, <span style="text-decoration: underline;">msofla</span>, <span style="text-decoration: underline;">msoiow</span>, <span style="text-decoration: underline;">msomin</span>, <span style="text-decoration: underline;">msoawx</span>, <span style="text-decoration: underline;">msonos</span>, <span style="text-decoration: underline;">msoapg</span>, <span style="text-decoration: underline;">msowfy</span>,&nbsp;<span style="text-decoration: underline;">msohad</span>, <span style="text-decoration: underline;">msoaws</span>, <span style="text-decoration: underline;">msoien</span>, <span style="text-decoration: underline;">msokla</span>, <span style="text-decoration: underline;">msocol</span>,&nbsp;<span style="text-decoration: underline;">msowtx</span>, <span style="text-decoration: underline;">msowis</span>, <span style="text-decoration: underline;">msolju</span>, <span style="text-decoration: underline;">mso470</span>, <span style="text-decoration: underline;">msodcn</span>, <span style="text-decoration: underline;">msoind</span>, <span style="text-decoration: underline;">msoflt</span>, <span style="text-decoration: underline;">msoalk</span>, <span style="text-decoration: underline;">msogeo</span>, <span style="text-decoration: underline;">msovir</span>, <span style="text-decoration: underline;">msomca</span>, <span style="text-decoration: underline;">msothr</span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">proflr</span><span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">prflr,
prflrb, prflrj<sup>1,3</sup>, prflrp</span><span style="font-family: Courier New;"></span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">qkscat</td>


















      <td style="font-family: Courier New; font-style: italic;">o</td>


















      <td style="font-family: Courier New; font-style: italic;">qscat</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">rassda<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R,N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">rass<br>


















      </td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">rtovs</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">o</td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic; color: rgb(0, 0, 0);">rtovs</td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">satwnd</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: courier new;"><span style="font-weight: bold;">R</span></span><sup><span style="font-size: 10pt;"><span style="font-family: courier new;"><span style="font-weight: bold;">8</span></span></span></sup><span style="font-family: courier new;"><sup><span style="font-weight: bold;"></span></sup>,<span style="font-weight: bold;">N</span></span><sup><span style="font-size: 10pt;"><span style="font-family: courier new;"><span style="font-weight: bold;">8</span></span></span></sup><span style="font-family: courier new;"><span style="font-weight: bold;"></span>,<span style="font-weight: bold;">G<sup>8</sup></span>,<span style="font-weight: bold;">F<sup>8</sup></span>,<span style="font-weight: bold;">C</span>,<span style="font-weight: bold;">M</span></span><sup><span style="font-size: 10pt;"><span style="font-family: courier new;"><span style="font-weight: bold;">8</span></span></span></sup></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">infus,
h2ius, visus, 3p9us<sup>12</sup>, infin</span><span style="font-family: Courier New;"><sup>1,3,11</sup>,
visin</span><span style="font-family: Courier New;"><sup>1,3,11</sup></span><span style="font-family: Courier New;">,
h20in</span><span style="font-family: Courier New;"><sup>1,3,11</sup></span><span style="font-family: Courier New;">,
infja</span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;">,
visja</span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;">,
h20ja</span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;">,
infeu</span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;">, viseu</span><sup><span style="font-size: 10pt;"><span style="font-family: Courier New;"></span></span></sup><span style="font-family: Courier New;">, h20eu</span><sup><span style="font-size: 10pt;"><span style="font-family: Courier New;"></span></span></sup><span style="font-family: Courier New;">, infmo, h20mo, infav<sup>12</sup>,
infvr<sup>12</sup>, infusr<sup>12</sup>,&nbsp;h2dusr<sup>12</sup>,&nbsp;visusr<sup>12</sup>,&nbsp;h2tusr<sup>12</sup>,&nbsp;3p9usr<sup>12</sup><br>


















      </span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;"></span><span style="font-family: Courier New;"></span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0); font-style: italic;"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">sfcbog</span><span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="color: rgb(0, 0, 0); font-style: italic;"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">slpbg</span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">sfcshp</span><span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">C</span>,<span style="font-weight: bold;">M</span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;"><span style="text-decoration: underline;">ships</span>,
shipsu, dbuoy, mbuoy, lcman, tideg, cstgd<sup>12</sup></span><span style="font-size: 10pt;"><span style="font-family: Courier New;"></span></span><span style="font-family: Courier New;"> </span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">ssmip</td>


















      <td style="font-family: Courier New; font-style: italic;">o</td>


















      <td style="font-family: Courier New; font-style: italic;">ssmip</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">ssmipn</td>


















      <td style="font-family: Courier New; font-style: italic;">o</td>


















      <td style="font-family: Courier New; font-style: italic;">ssmipn</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">ssmit</td>


















      <td style="font-family: Courier New; font-style: italic;">o</td>


















      <td style="font-family: Courier New; font-style: italic;">ssmit</td>


















    </tr>


















    <tr valign="top">


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">vadwnd</span><span style="font-size: 10pt;"></span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: courier new;"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</span></td>


















      <td style="color: rgb(0, 0, 0);"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">nxrdw,&nbsp;nxrdw2</span><sup><span style="font-size: 10pt;"><span style="font-family: Courier New;">2,5</span></span></sup><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="color: rgb(0, 0, 0); font-family: Courier New; font-style: italic;">wndsat</td>


















      <td style="color: rgb(0, 0, 0); font-family: Courier New; font-style: italic;"><span style="font-weight: bold;"></span><sup><span style="font-size: 10pt;"><span style="font-size: 10pt; font-weight: bold;"></span></span></sup><span style="font-weight: bold;"></span><sup><span style="font-size: 10pt; font-weight: bold;"></span></sup><span style="font-weight: bold;"></span><span style="font-weight: bold;"></span><span style="font-weight: bold;"></span></td>


















      <td style="color: rgb(0, 0, 0); font-family: Courier New; font-style: italic;">wdsat</td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















</p>


















</span><span style="font-size: 10pt;">
<p><span style="font-size: 10pt;"></span><br>


















</p>


















<hr width="100%"><br>


















<a name="c"></a><br>


















&nbsp;
</span></p>


















<p style="font-family: courier new;"><big><span style="font-family: times new roman;">Table 1.c&nbsp;&nbsp; Data group
mnemonics used to generate BUFR
dump
files in the various NCEP networks.&nbsp; These dump files are then
read
by the subsequent analysis codes (with the exception of "satwnd", they
do not pass through the PREPBUFR
processing steps) (last revised 2/11/2018 <span style="font-style: italic;">- not completely up to date!</span>).</span>
</big><br>


















&nbsp;
</p>


















<p style="font-family: courier new;">Key for NETWORK ("NET") column -
if&nbsp;<span style="font-weight: bold;">BOLDFACE AND UPPER-CASE&nbsp;</span>indicates
the dump file for this group is read in by the
subsequent
analysis
codes and at least some data in the dump file is actually assimilated
(not just monitored) by the analysis; if <span style="font-style: italic;">italics</span>&nbsp;indicates
the dump file for this group is normally dumped in this network but is
temporarily not available (in this case may also be in <span style="font-style: italic;">italics</span> in either "GROUP MENMONIC"
or&nbsp;"MNEMONICS INCLUDED" columns or both):
<br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-weight: bold;">C</span>/c -
group is
dumped in CDAS network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-weight: bold;">F</span>/f -
group is
dumped in GDAS&nbsp;network<br>


















&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-weight: bold;">G</span>/g -
group is
dumped in GFS&nbsp;network<br>


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp; M/m -
group is dumped in RTMA and&nbsp;URMA networks<br>


















</span>&nbsp;&nbsp;&nbsp;&nbsp; <span style="font-weight: bold;">N</span>/n
-
group is
dumped in NAM&nbsp;network<br>


















<span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;</span><span style="font-style: italic; font-family: courier new;">o &nbsp; - group
is
obsolete and is not dumped in any network (also in italics)</span><br>


















<span style="font-family: courier new;">&nbsp; &nbsp;&nbsp; <span style="font-weight: bold;">R</span>/r -
group is dumped in&nbsp;RAP network (all runs except </span><span style="font-family: courier new;">Early-cycle-HRRR)</span><br>













<span style="font-family: courier new;">&nbsp; &nbsp; &nbsp;<span style="font-weight: bold;">H</span>/r - </span><span style="font-family: courier new;">group is dumped in&nbsp;RAP Early-cycle-HRRR run<br>













</span>&nbsp;&nbsp;&nbsp;&nbsp;&nbsp;<span style="font-weight: bold;"></span><span style="font-style: italic;">t
&nbsp; - group
consists
of future data types and is currently not dumped in any network (also
in
italics)</span><br>


















</p>


















<span style="font-family: courier new;"><br>


















Key for superscripts in "NET" column:</span><a style="font-family: courier new;" name="c.2"></a><span style="font-family: courier new;"><br>


















&nbsp; &nbsp;&nbsp; 1 - input to
TRMM TMI reprocessing program BUFR_SUPERTMI which outputs superobed
data
(on a 1 degree lat/lon grid) in a file called "sptrmm&rdquo; which is
read by
the subsequent analysis codes if network is <span style="font-weight: bold;">boldface</span><span style="font-weight: bold;"></span><br>


















<br>


















<br>


















Key for superscripts in "MNEMONICS INCLUDED" column:<br>


















&nbsp;&nbsp;&nbsp;&nbsp; 1 - only included if reports are within the
selected dump time window<br>


















</span><span style="font-family: courier new;">&nbsp; &nbsp; &nbsp;2 -
not included in&nbsp;RAP network dumps<br>


















</span><span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;&nbsp;
3 -
not included in NAM&nbsp;network dumps<br>


















</span><span style="font-family: courier new;">&nbsp;&nbsp;&nbsp;
&nbsp;4 -
not included in RTMA and&nbsp;URMA network dumps<br>















&nbsp; &nbsp; &nbsp;5 - included only in GFS and GDAS network dumps<br>


















</span><span style="font-size: 10pt;">
<p>&nbsp;&nbsp;
<br>


















&nbsp;
<table style="width: 100%;" border="1">


















  <tbody>


















    <tr valign="top">


















      <td><span style="font-size: 10pt;"></span><span style="font-size: 10pt;"></span><span style="font-size: 10pt;">GROUP
MNEMONIC</span> <br>


















      <span style="font-size: 10pt;">(dump file)</span></td>


















      <td><span style="font-size: 10pt;">NET</span></td>


















      <td><span style="font-size: 10pt;">MNEMONICS INCLUDED</span><span style="font-size: 10pt;"><span style="font-size: 10pt;"> (<span style="text-decoration: underline;">underlined</span> means some or
all reports in this mnemonic&nbsp;are <a href="http://www.nco.ncep.noaa.gov/sib/restricted_data/restricted_data_pmb/">restricted
with respect to redistribution outside of NCEP for some amount of time</a>)</span></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">airsev</td>


















      <td style="font-family: Courier New;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">airsev</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">amsr2</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">amsr2</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">amsre<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">g,f,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; font-style: italic;">amsre<br>


















      </td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">atms</td>


















      <td style="font-family: Courier New;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">atms</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">atmsdb</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">atmsdb</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;" align="left" valign="top">avcsam</td>


















      <td style="font-family: Courier New;" align="left" valign="top">g,f,c</td>


















      <td style="font-family: Courier New;" align="left" valign="top">avcsam</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;" align="left" valign="top">avcspm</td>


















      <td style="font-family: Courier New;" align="left" valign="top">g,f,c</td>


















      <td style="font-family: Courier New;" align="left" valign="top">avcspm</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">bathy</td>


















      <td style="font-family: Courier New;">g,f,c</td>


















      <td style="font-family: Courier New;">bathy</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">cris</td>


















      <td style="font-family: Courier New;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">cris</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">crisdb</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">crisdb</td>


















    </tr>


















    <tr>















      <td><span style="font-family: Courier New;">crisf4</span></td>















      <td style="font-family: Courier New;">g,f</td>















      <td style="font-family: Courier New;">crisf4</td>















    </tr>















    <tr>


















      <td style="font-family: Courier New;">efclam</td>


















      <td style="font-family: Courier New;"><span style="font-weight: bold;">M</span></td>


















      <td style="font-family: Courier New;">efclam</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">esamua</td>


















      <td style="font-family: Courier New;">r,n,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">esamua</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">esatms</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">esatms</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">escris</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">escris</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">eshrs3</td>


















      <td style="font-family: Courier New;">r,n,g,f,c</td>


















      <td style="font-family: Courier New;">eshrs3</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">esiasi</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">esiasi</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">esmhs</td>


















      <td style="font-family: Courier New;">r,n,g,f,c</td>


















      <td style="font-family: Courier New;">esmhs</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new;">geoimr<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);">g,f,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new;">geoimr<br>


















      </td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">goesfv</td>


















      <td style="font-family: Courier New;"><span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">geost1</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;" align="left" valign="top">gome</td>


















      <td style="font-family: Courier New;" align="left" valign="top">g,f,c</td>


















      <td style="font-family: Courier New;" align="left" valign="top">gome</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">gpsro</td>


















      <td style="font-family: Courier New;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">gpsro</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">iasidb</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">iasidb</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">lghtng</td>


















      <td style="font-family: Courier New;"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,c</td>


















      <td style="font-family: Courier New;">ltngsr,&nbsp;ltnglr</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">lgycld</td>


















      <td style="font-family: Courier New;"><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,c</td>


















      <td style="font-family: Courier New;">lgycld</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; font-style: italic;">mls</td>


















      <td style="font-family: Courier New; font-style: italic;">g,f,c</td>


















      <td style="font-family: Courier New; font-style: italic;">mls
&nbsp;<span style="font-weight: bold; color: rgb(255, 0, 0);">--&gt;
empty as of 12z 01/31/2017, no longer even dumped after 02/10/2017</span></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;" align="left" valign="top">mtiasi</td>


















      <td style="font-family: Courier New;" align="left" valign="top"><span style="font-size: 10pt;">r,</span><span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;" align="left" valign="top">mtiasi</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new; height: 133px;">nexrad<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; height: 133px;"><span style="font-weight: bold;">H</span>,<span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new; height: 133px;">rd2w00<sup><span style="font-size: 10pt;">1</span></sup>,
rd2w01<span style="font-size: 10pt;"><span style="font-size: 10pt;"></span></span><sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w02<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w03<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w04<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w05<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w06<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w07<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w08<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w09<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w10<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w11<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w12<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w13<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w14<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w15<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w16<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w17<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w18<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w19<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w20<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w21<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w22<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2w23<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1</span></span></sup>,
rd2r00<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r01<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r02<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r03<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r04<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r05<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r06<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r07<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r08<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r09<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r10<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r11<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r12<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r13<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r14<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r15<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r16<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r17<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r18<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r19<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r20<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r21<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r22<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>,
rd2r23<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;">1,2</span></span></sup>
      </td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">omi</td>


















      <td style="font-family: Courier New;"><span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">omi</td>


















    </tr>


















    <tr valign="top">


















      <td style="font-family: courier new; font-style: italic;">osbuv</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="font-family: courier new; font-style: italic;">osbuv</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">osbuv8</td>


















      <td style="font-family: Courier New;">r,n,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">osbuv8</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new;">radwnd</td>


















      <td style="vertical-align: top; font-family: courier new; color: rgb(0, 0, 0);"><span style="font-weight: bold;"></span><span style="font-weight: bold;"></span>r,n,c</td>


















      <td style="vertical-align: top; font-family: courier new;">radw30,
radw25</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">saphir</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">saphir</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New; vertical-align: top;">satwnd</td>


















      <td style="font-family: Courier New; vertical-align: top;"><span style="font-weight: bold;"></span><span style="font-weight: bold;">R</span>,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,<span style="font-weight: bold;">M</span><span style="font-size: 10pt;"><sup><span style="font-size: 10pt;"><span style="font-family: courier new;"><span style="font-weight: bold;"></span></span></span></sup></span></td>


















      <td style="font-family: Courier New; vertical-align: top;">infus,
h2ius, visus, 3p9us, infin<sup><span style="font-family: courier new;">2,3,4</span></sup>,
visin<sup><span style="font-family: courier new;">2,3,4</span></sup>,
h20in<sup><span style="font-family: courier new;">2,3,4</span></sup>,
infja, visja, h20ja, infeu, viseu,
h20eu, infmo, h20mo, infav, infvr, infusr<sup><sub><span style="font-size: 10pt;"><span style="font-family: courier new;">5</span></span></sub></sup>,&nbsp;h2dusr<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-family: courier new;">5</span></span></span></sup>,&nbsp;visusr<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-family: courier new;">5</span></span></span></sup>,&nbsp;h2tusr<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-family: courier new;">5</span></span></span></sup>,&nbsp;3p9usr<sup><span style="font-size: 10pt;"><span style="font-size: 10pt;"><span style="font-family: courier new;">5</span></span></span></sup></td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">sevasr</td>


















      <td style="font-family: Courier New;">g,f</td>


















      <td style="font-family: Courier New;">sevasr</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">sevcsr</td>


















      <td style="font-family: Courier New;">r<span style="font-weight: bold;">,N,G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">sevcsr</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">ssmisu</td>


















      <td style="font-family: Courier New;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: Courier New;">ssmisu</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">tesac</td>


















      <td style="font-family: Courier New;">g,f,c</td>


















      <td style="font-family: Courier New;">tesac</td>


















    </tr>


















    <tr>


















      <td style="font-family: Courier New;">trkob</td>


















      <td style="font-family: Courier New;">g,f,c</td>


















      <td style="font-family: Courier New;">trkob</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; height: 24px; font-style: italic;">trmm</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); height: 24px; font-style: italic;"><span style="font-weight: bold;">o</span><sup></sup></td>


















      <td style="font-family: courier new; height: 24px; font-style: italic;">trmm</td>


















    </tr>


















    <tr valign="top">


















      <td style="font-style: italic;"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">1bhrs2</span><span style="font-size: 10pt;"></span></td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="font-style: italic;"><span style="font-size: 10pt;"></span><span style="font-family: Courier New;">1bhrs2</span><span style="font-size: 10pt;"></span></td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic;">1bmsu</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="font-family: courier new; font-style: italic;">1bmsu</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new;">1bamua</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0);">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c</td>


















      <td style="font-family: courier new;">1bamua</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic;">1bamub</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="font-family: courier new; font-style: italic;">1bamub</td>


















    </tr>


















    <tr>


















      <td style="font-family: courier new; font-style: italic;">1bhrs3</td>


















      <td style="font-family: courier new; color: rgb(0, 0, 0); font-style: italic;">o</td>


















      <td style="font-family: courier new; font-style: italic;">1bhrs3</td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new;">1bhrs4<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new;">r,n,g,f,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new;">1bhrs4<br>


















      </td>


















    </tr>


















    <tr>


















      <td style="vertical-align: top; font-family: courier new;">1bmhs<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new;">r,<span style="font-weight: bold;">N</span>,<span style="font-weight: bold;">G</span>,<span style="font-weight: bold;">F</span>,c<br>


















      </td>


















      <td style="vertical-align: top; font-family: courier new;">1bmhs<br>


















      </td>


















    </tr>


















  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  </tbody>
</table>


















<br>


















&nbsp;
<br>


















</p>


















</span>
<br>


















<br>


















</body>
</html>
